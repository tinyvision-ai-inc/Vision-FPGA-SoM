`timescale 1ps/1ps
module RAM40_16KNR ( RDATA, RCLKN, RCLKE, RE, RADDR, WCLK, WCLKE, WE, WADDR, MASK, WDATA ); 

output	[15:0]	RDATA;  
input         	RCLKN;   
input           RCLKE; 
input           RE; 
input	[12:0]  RADDR; 
input           WCLK; 
input           WCLKE; 
input           WE; 
input 	[12:0]  WADDR; 
input 	[15:0]  MASK; 
input 	[15:0]	WDATA; 

parameter WRITE_MODE = 0;    // Configure Write Port as 1024x16 (0)/ 20148x8 (1)/ 4096x4 (2)/ 8192x2 (3)     
parameter READ_MODE  = 0;    // Configure Read  Port as 1024x16 (0)/ 20148x8 (1)/ 4096x4 (2)/ 8192x2 (3)

parameter INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;


wire RCLK;
assign (weak0, weak1) RCLKE =1'b1 ;
assign (weak0, weak1) RE =1'b0 ;
assign (weak0, weak1) WCLKE =1'b1 ;
assign (weak0, weak1) WE =1'b0 ;
assign RCLK = ~RCLKN;

RAM40_16K ram40mh_16K_nr_inst (
	.RDATA(RDATA),
	.RCLK(RCLK),
	.RCLKE(RCLKE),
	.RE(RE),
	.RADDR(RADDR),
	.WCLK(WCLK),
	.WCLKE(WCLKE),
	.WE(WE),
	.WADDR(WADDR),
	.MASK(MASK),
	.WDATA(WDATA));

defparam ram40mh_16K_nr_inst.WRITE_MODE = WRITE_MODE;
defparam ram40mh_16K_nr_inst.READ_MODE = READ_MODE;

defparam ram40mh_16K_nr_inst.INIT_0 = INIT_0;
defparam ram40mh_16K_nr_inst.INIT_1 = INIT_1;
defparam ram40mh_16K_nr_inst.INIT_2 = INIT_2;
defparam ram40mh_16K_nr_inst.INIT_3 = INIT_3;
defparam ram40mh_16K_nr_inst.INIT_4 = INIT_4;
defparam ram40mh_16K_nr_inst.INIT_5 = INIT_5;
defparam ram40mh_16K_nr_inst.INIT_6 = INIT_6;
defparam ram40mh_16K_nr_inst.INIT_7 = INIT_7;
defparam ram40mh_16K_nr_inst.INIT_8 = INIT_8;
defparam ram40mh_16K_nr_inst.INIT_9 = INIT_9;
defparam ram40mh_16K_nr_inst.INIT_A = INIT_A;
defparam ram40mh_16K_nr_inst.INIT_B = INIT_B;
defparam ram40mh_16K_nr_inst.INIT_C = INIT_C;
defparam ram40mh_16K_nr_inst.INIT_D = INIT_D;
defparam ram40mh_16K_nr_inst.INIT_E = INIT_E;
defparam ram40mh_16K_nr_inst.INIT_F = INIT_F;

defparam ram40mh_16K_nr_inst.INIT_0 = INIT_0;
defparam ram40mh_16K_nr_inst.INIT_1 = INIT_1;
defparam ram40mh_16K_nr_inst.INIT_2 = INIT_2;
defparam ram40mh_16K_nr_inst.INIT_3 = INIT_3;
defparam ram40mh_16K_nr_inst.INIT_4 = INIT_4;
defparam ram40mh_16K_nr_inst.INIT_5 = INIT_5;
defparam ram40mh_16K_nr_inst.INIT_6 = INIT_6;
defparam ram40mh_16K_nr_inst.INIT_7 = INIT_7;
defparam ram40mh_16K_nr_inst.INIT_8 = INIT_8;
defparam ram40mh_16K_nr_inst.INIT_9 = INIT_9;
defparam ram40mh_16K_nr_inst.INIT_A = INIT_A;
defparam ram40mh_16K_nr_inst.INIT_B = INIT_B;
defparam ram40mh_16K_nr_inst.INIT_C = INIT_C;
defparam ram40mh_16K_nr_inst.INIT_D = INIT_D;
defparam ram40mh_16K_nr_inst.INIT_E = INIT_E;
defparam ram40mh_16K_nr_inst.INIT_F = INIT_F;

defparam ram40mh_16K_nr_inst.INIT_0 = INIT_0;
defparam ram40mh_16K_nr_inst.INIT_1 = INIT_1;
defparam ram40mh_16K_nr_inst.INIT_2 = INIT_2;
defparam ram40mh_16K_nr_inst.INIT_3 = INIT_3;
defparam ram40mh_16K_nr_inst.INIT_4 = INIT_4;
defparam ram40mh_16K_nr_inst.INIT_5 = INIT_5;
defparam ram40mh_16K_nr_inst.INIT_6 = INIT_6;
defparam ram40mh_16K_nr_inst.INIT_7 = INIT_7;
defparam ram40mh_16K_nr_inst.INIT_8 = INIT_8;
defparam ram40mh_16K_nr_inst.INIT_9 = INIT_9;
defparam ram40mh_16K_nr_inst.INIT_A = INIT_A;
defparam ram40mh_16K_nr_inst.INIT_B = INIT_B;
defparam ram40mh_16K_nr_inst.INIT_C = INIT_C;
defparam ram40mh_16K_nr_inst.INIT_D = INIT_D;
defparam ram40mh_16K_nr_inst.INIT_E = INIT_E;
defparam ram40mh_16K_nr_inst.INIT_F = INIT_F;

defparam ram40mh_16K_nr_inst.INIT_0 = INIT_0;
defparam ram40mh_16K_nr_inst.INIT_1 = INIT_1;
defparam ram40mh_16K_nr_inst.INIT_2 = INIT_2;
defparam ram40mh_16K_nr_inst.INIT_3 = INIT_3;
defparam ram40mh_16K_nr_inst.INIT_4 = INIT_4;
defparam ram40mh_16K_nr_inst.INIT_5 = INIT_5;
defparam ram40mh_16K_nr_inst.INIT_6 = INIT_6;
defparam ram40mh_16K_nr_inst.INIT_7 = INIT_7;
defparam ram40mh_16K_nr_inst.INIT_8 = INIT_8;
defparam ram40mh_16K_nr_inst.INIT_9 = INIT_9;
defparam ram40mh_16K_nr_inst.INIT_A = INIT_A;
defparam ram40mh_16K_nr_inst.INIT_B = INIT_B;
defparam ram40mh_16K_nr_inst.INIT_C = INIT_C;
defparam ram40mh_16K_nr_inst.INIT_D = INIT_D;
defparam ram40mh_16K_nr_inst.INIT_E = INIT_E;
defparam ram40mh_16K_nr_inst.INIT_F = INIT_F;

 
endmodule  // RAM40_16KNR 
