`timescale 10ps/1ps
module ClkMux (I, O);
input I;
output O;

	assign O = I;


endmodule
