`timescale 1ps/1ps
module LEDDA_IP ( LEDDCS,LEDDCLK,LEDDDAT7,LEDDDAT6,LEDDDAT5,LEDDDAT4,
	LEDDDAT3,LEDDDAT2,LEDDDAT1,LEDDDAT0,LEDDADDR3,LEDDADDR2,LEDDADDR1,
	LEDDADDR0,LEDDDEN,LEDDEXE,LEDDRST,PWMOUT0,PWMOUT1,PWMOUT2,LEDDON);	 
	
	input 	LEDDCS,LEDDCLK,LEDDDAT7,LEDDDAT6,LEDDDAT5,LEDDDAT4,LEDDDAT3,LEDDDAT2,
			LEDDDAT1,LEDDDAT0,LEDDADDR3,LEDDADDR2,LEDDADDR1,LEDDADDR0,LEDDDEN,LEDDEXE,LEDDRST; 
	output  PWMOUT0,PWMOUT1,PWMOUT2,LEDDON;
	
	wire LEDDCS, LEDDCLK,LEDDDAT7,LEDDDAT6,LEDDDAT5,LEDDDAT4,LEDDDAT3,LEDDDAT2, LEDDDAT1,LEDDDAT0,LEDDADDR3,LEDDADDR2,LEDDADDR1,LEDDADDR0,LEDDDEN,LEDDEXE,LEDDRST; 
	wire PWMOUT0,PWMOUT1,PWMOUT2,LEDDON;
	wire [7:0]  sb_ledd_dat={LEDDDAT7,LEDDDAT6,LEDDDAT5, LEDDDAT4,LEDDDAT3,LEDDDAT2,LEDDDAT1,LEDDDAT0};
	wire [3:0]	sb_ledd_adr={LEDDADDR3,LEDDADDR2,LEDDADDR1,LEDDADDR0};
	reg NOTIFIER;
	reg ledd_rst_async;
	initial
begin
   ledd_rst_async = 1'b1;
#100
   ledd_rst_async = 1'b0;
end
	ledd_ip_sub  ledd_ip_inst
	(
	.pwm_out_r(PWMOUT0),
	.pwm_out_g(PWMOUT1), 
	.pwm_out_b(PWMOUT2), 
	.ledd_on(LEDDON),
	.ledd_rst_async(ledd_rst_async), 
	.ledd_clk(LEDDCLK), 
	.ledd_cs(LEDDCS), 
	.ledd_den(LEDDDEN), 
	.ledd_adr(sb_ledd_adr), 
	.ledd_dat(sb_ledd_dat),
    .ledd_exe(LEDDEXE)
   );
   

   
endmodule
