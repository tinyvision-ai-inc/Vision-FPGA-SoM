`timescale 10ps/1ps
module CascadeBuf(I, O);
input I;
output O;

assign O = I;


endmodule
