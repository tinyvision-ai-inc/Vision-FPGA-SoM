`timescale 1ns/1ns
module VLO ( Z );
    output Z ;
  supply0 VSS;
  buf (Z , VSS);
endmodule
