`timescale 10ps/1ps
module IpInMux(I, O);
input I;
output O;

assign O = I;


endmodule
