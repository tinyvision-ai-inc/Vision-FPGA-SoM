`timescale 10ps/1ps
module Glb2LocalMux(I, O);
input I;
output O;

	assign O = I;
	

endmodule
