`timescale 10ps/1ps
module GlobalMux(I, O);
input I;
output O;

	assign O = I;


endmodule
