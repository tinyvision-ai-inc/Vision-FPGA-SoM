`timescale 1ps/1ps
module ICE_IR500_DRV   (
	IRLEDEN,
	IRPWM,
	CURREN,
	IRLEDEN2,
	IRPWM2,
	IRLED1,
	IRLED2
);

parameter IR500_CURRENT = "0b000000000000";
parameter CURRENT_MODE = "0b0";

	input IRLEDEN;
	input IRPWM;
	input CURREN;
	input IRLEDEN2;
	input IRPWM2;
	output IRLED1;
	output IRLED2;

 ICE_IR500_DRV_CORE #(.IR500_CURRENT(IR500_CURRENT),.CURRENT_MODE(CURRENT_MODE))
inst
 (
	.CURREN(CURREN),
	.IRLEDEN(IRLEDEN),
	.IRPWM(IRPWM),
	.IRLEDEN2(IRLEDEN2),
	.IRPWM2(IRPWM2),
	.IRLED1(IRLED1),
	.IRLED2(IRLED2)
);
endmodule
