`timescale 10ps/1ps
module Span4Mux(I, O);
input I;
output O;

	assign O = I;
	

endmodule
