`timescale 10ps/1ps
module ColCtrlBuf(I, O);
input I;
output O;

	assign O = I;


endmodule
