`timescale 10ps/1ps
module InMux(I, O);
input I;
output O;

	assign O = I;

endmodule
