`timescale 10ps/1ps
module G2TBuf (I, O);
parameter X = 1;
parameter Y = 1;
input I;
output O;
   assign O = I ;


endmodule
