`timescale 1ns/1ns
module VFB_B (ADDRESS13, ADDRESS12, ADDRESS11, ADDRESS10, ADDRESS9, ADDRESS8, ADDRESS7, ADDRESS6, ADDRESS5, ADDRESS4, ADDRESS3, ADDRESS2, ADDRESS1, ADDRESS0, DATAIN15, DATAIN14, DATAIN13, DATAIN12, DATAIN11, DATAIN10, DATAIN9, DATAIN8, DATAIN7, DATAIN6, DATAIN5, DATAIN4, DATAIN3, DATAIN2, DATAIN1, DATAIN0, MASKWREN3, MASKWREN2, MASKWREN1, MASKWREN0, WREN, CHIPSELECT, CLOCK, RDMARGINEN, RDMARGIN3, RDMARGIN2, RDMARGIN1, RDMARGIN0, STANDBY, SLEEP, POWEROFF_N, TEST, DATAOUT15, DATAOUT14, DATAOUT13, DATAOUT12, DATAOUT11, DATAOUT10, DATAOUT9, DATAOUT8, DATAOUT7, DATAOUT6, DATAOUT5, DATAOUT4, DATAOUT3, DATAOUT2, DATAOUT1, DATAOUT0);

	//Port Type List [Expanded Bus/Bit]
	input ADDRESS13;
	input ADDRESS12;
	input ADDRESS11;
	input ADDRESS10;
	input ADDRESS9;
	input ADDRESS8;
	input ADDRESS7;
	input ADDRESS6;
	input ADDRESS5;
	input ADDRESS4;
	input ADDRESS3;
	input ADDRESS2;
	input ADDRESS1;
	input ADDRESS0;
	input DATAIN15;
	input DATAIN14;
	input DATAIN13;
	input DATAIN12;
	input DATAIN11;
	input DATAIN10;
	input DATAIN9;
	input DATAIN8;
	input DATAIN7;
	input DATAIN6;
	input DATAIN5;
	input DATAIN4;
	input DATAIN3;
	input DATAIN2;
	input DATAIN1;
	input DATAIN0;
	input MASKWREN3;
	input MASKWREN2;
	input MASKWREN1;
	input MASKWREN0;
	input WREN;
	input CHIPSELECT;
	input CLOCK;
	input RDMARGINEN;
	input RDMARGIN3;
	input RDMARGIN2;
	input RDMARGIN1;
	input RDMARGIN0;
	input STANDBY;
	input SLEEP;
	input POWEROFF_N;
	input TEST;
	output DATAOUT15;
	output DATAOUT14;
	output DATAOUT13;
	output DATAOUT12;
	output DATAOUT11;
	output DATAOUT10;
	output DATAOUT9;
	output DATAOUT8;
	output DATAOUT7;
	output DATAOUT6;
	output DATAOUT5;
	output DATAOUT4;
	output DATAOUT3;
	output DATAOUT2;
	output DATAOUT1;
	output DATAOUT0;


	//Assigning input IP Ports to corresponding SW bit ports [Inputs]
	wire [13:0] ADDRESS;
	assign ADDRESS = {ADDRESS13, ADDRESS12, ADDRESS11, ADDRESS10, ADDRESS9, ADDRESS8, ADDRESS7, ADDRESS6, ADDRESS5, ADDRESS4, ADDRESS3, ADDRESS2, ADDRESS1, ADDRESS0};
	wire [15:0] DATAIN;
	assign DATAIN = {DATAIN15, DATAIN14, DATAIN13, DATAIN12, DATAIN11, DATAIN10, DATAIN9, DATAIN8, DATAIN7, DATAIN6, DATAIN5, DATAIN4, DATAIN3, DATAIN2, DATAIN1, DATAIN0};
	wire [3:0] MASKWREN;
	assign MASKWREN = {MASKWREN3, MASKWREN2, MASKWREN1, MASKWREN0};
	wire [3:0] RDMARGIN;
	assign RDMARGIN = {RDMARGIN3, RDMARGIN2, RDMARGIN1, RDMARGIN0};
	//Fanning IP Bus Output to Individual SW Bit [Outputs]
	wire [15:0] DATAOUT;
	assign DATAOUT0 = DATAOUT[0];
	assign DATAOUT1 = DATAOUT[1];
	assign DATAOUT2 = DATAOUT[2];
	assign DATAOUT3 = DATAOUT[3];
	assign DATAOUT4 = DATAOUT[4];
	assign DATAOUT5 = DATAOUT[5];
	assign DATAOUT6 = DATAOUT[6];
	assign DATAOUT7 = DATAOUT[7];
	assign DATAOUT8 = DATAOUT[8];
	assign DATAOUT9 = DATAOUT[9];
	assign DATAOUT10 = DATAOUT[10];
	assign DATAOUT11 = DATAOUT[11];
	assign DATAOUT12 = DATAOUT[12];
	assign DATAOUT13 = DATAOUT[13];
	assign DATAOUT14 = DATAOUT[14];
	assign DATAOUT15 = DATAOUT[15];

	//IP Ports Tied Off for Simulation
	//Attribute List
	`include "convertDeviceString.v"

	SPRAM256KA SRAM_inst(.ADDRESS(ADDRESS), .DATAIN(DATAIN), .MASKWREN(MASKWREN), .WREN(WREN), .CHIPSELECT(CHIPSELECT), .CLOCK(CLOCK), .RDMARGINEN(RDMARGINEN), .RDMARGIN(RDMARGIN), .STANDBY(STANDBY), .SLEEP(SLEEP), .POWEROFF(POWEROFF_N), .TEST(TEST), .DATAOUT(DATAOUT));


endmodule
