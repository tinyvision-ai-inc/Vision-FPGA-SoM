`timescale 10ps/1ps
module IoSpan4Mux(I, O);
input I;
output O;

	assign O = I;
	

endmodule
