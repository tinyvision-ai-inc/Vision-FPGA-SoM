`timescale 10ps/1ps
module Span12Mux_s10_v(I, O);
input I;
output O;

	assign O = I;
	

endmodule
