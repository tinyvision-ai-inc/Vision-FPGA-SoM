`timescale 1ps/1ps
module WARMBOOT_SUB (	
BOOT, S1, S0);

input BOOT;
input S1;
input S0;			

endmodule	//WARMBOOT_SUB
