`timescale 10ps/1ps
module Span12Mux_s3_h(I, O);
input I;
output O;

	assign O = I;
	

endmodule
