`timescale 10ps/1ps
module gio2CtrlBuf(I, O);
input I;
output O;

	assign O = I;


endmodule
