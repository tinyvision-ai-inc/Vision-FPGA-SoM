`timescale 1ns/1ns
module PLL_B (REFERENCECLK, FEEDBACK, DYNAMICDELAY7, DYNAMICDELAY6, DYNAMICDELAY5, DYNAMICDELAY4, DYNAMICDELAY3, DYNAMICDELAY2, DYNAMICDELAY1, DYNAMICDELAY0, BYPASS, RESET_N, SCLK, SDI, LATCH, INTFBOUT, OUTCORE, OUTGLOBAL, OUTCOREB, OUTGLOBALB, SDO, LOCK);

	//Port Type List [Expanded Bus/Bit]
	input REFERENCECLK;
	input FEEDBACK;
	input DYNAMICDELAY7;
	input DYNAMICDELAY6;
	input DYNAMICDELAY5;
	input DYNAMICDELAY4;
	input DYNAMICDELAY3;
	input DYNAMICDELAY2;
	input DYNAMICDELAY1;
	input DYNAMICDELAY0;
	input BYPASS;
	input RESET_N;
	input SCLK;
	input SDI;
	input LATCH;
	output INTFBOUT;
	output OUTCORE;
	output OUTGLOBAL;
	output OUTCOREB;
	output OUTGLOBALB;
	output SDO;
	output LOCK;


	//Assigning input IP Ports to corresponding SW bit ports [Inputs]
	wire [7:0] DYNAMICDELAY;
	assign DYNAMICDELAY = {DYNAMICDELAY7, DYNAMICDELAY6, DYNAMICDELAY5, DYNAMICDELAY4, DYNAMICDELAY3, DYNAMICDELAY2, DYNAMICDELAY1, DYNAMICDELAY0};

	//IP Ports Tied Off for Simulation
	//Attribute List
	parameter FEEDBACK_PATH = "SIMPLE";
	parameter DELAY_ADJUSTMENT_MODE_FEEDBACK = "FIXED";
	parameter FDA_FEEDBACK = "0";
	parameter DELAY_ADJUSTMENT_MODE_RELATIVE = "FIXED";
	parameter FDA_RELATIVE = "0";
	parameter SHIFTREG_DIV_MODE = "0";
	parameter PLLOUT_SELECT_PORTA = "SHIFTREG_0deg";
	parameter PLLOUT_SELECT_PORTB = "SHIFTREG_0deg";
	parameter DIVR = "0";
	parameter DIVF = "0";
	parameter DIVQ = "1";
	parameter FILTER_RANGE = "0";
	parameter EXTERNAL_DIVIDE_FACTOR = "NONE";
	parameter ENABLE_ICEGATE_PORTA = "0";
	parameter ENABLE_ICEGATE_PORTB = "0";
	parameter TEST_MODE = "0";
	parameter FREQUENCY_PIN_REFERENCECLK = "NONE";
	`include "convertDeviceString.v"
	//Converted Attribute List [For Device Binary / Hex String]
	localparam CONVERTED_FDA_FEEDBACK = convertDeviceString(FDA_FEEDBACK);
	localparam CONVERTED_FDA_RELATIVE = convertDeviceString(FDA_RELATIVE);
	localparam CONVERTED_SHIFTREG_DIV_MODE = convertDeviceString(SHIFTREG_DIV_MODE);
	localparam CONVERTED_DIVR = convertDeviceString(DIVR);
	localparam CONVERTED_DIVF = convertDeviceString(DIVF);
	localparam CONVERTED_DIVQ = convertDeviceString(DIVQ);
	localparam CONVERTED_FILTER_RANGE = convertDeviceString(FILTER_RANGE);
	localparam CONVERTED_ENABLE_ICEGATE_PORTA = convertDeviceString(ENABLE_ICEGATE_PORTA);
	localparam CONVERTED_ENABLE_ICEGATE_PORTB = convertDeviceString(ENABLE_ICEGATE_PORTB);
	localparam CONVERTED_TEST_MODE = convertDeviceString(TEST_MODE);

	PLL40_2F_CORE PLL_inst(.REFERENCECLK(REFERENCECLK), .EXTFEEDBACK(FEEDBACK), .DYNAMICDELAY(DYNAMICDELAY), .BYPASS(BYPASS), .RESETB(RESET_N), .SCLK(SCLK), .SDI(SDI), .LATCHINPUTVALUE(LATCH), .PLLOUTCOREA(OUTCORE), .PLLOUTGLOBALA(OUTGLOBAL), .PLLOUTCOREB(OUTCOREB), .PLLOUTGLOBALB(OUTGLOBALB), .SDO(SDO), .LOCK(LOCK));
	defparam PLL_inst.FEEDBACK_PATH = FEEDBACK_PATH;
	defparam PLL_inst.DELAY_ADJUSTMENT_MODE_FEEDBACK = DELAY_ADJUSTMENT_MODE_FEEDBACK;
	defparam PLL_inst.FDA_FEEDBACK = CONVERTED_FDA_FEEDBACK;
	defparam PLL_inst.DELAY_ADJUSTMENT_MODE_RELATIVE = DELAY_ADJUSTMENT_MODE_RELATIVE;
	defparam PLL_inst.FDA_RELATIVE = CONVERTED_FDA_RELATIVE;
	defparam PLL_inst.SHIFTREG_DIV_MODE = CONVERTED_SHIFTREG_DIV_MODE;
	defparam PLL_inst.PLLOUT_SELECT_PORTA = PLLOUT_SELECT_PORTA;
	defparam PLL_inst.PLLOUT_SELECT_PORTB = PLLOUT_SELECT_PORTB;
	defparam PLL_inst.DIVR = CONVERTED_DIVR;
	defparam PLL_inst.DIVF = CONVERTED_DIVF;
	defparam PLL_inst.DIVQ = CONVERTED_DIVQ;
	defparam PLL_inst.FILTER_RANGE = CONVERTED_FILTER_RANGE;
	defparam PLL_inst.EXTERNAL_DIVIDE_FACTOR = EXTERNAL_DIVIDE_FACTOR;
	defparam PLL_inst.ENABLE_ICEGATE_PORTA = CONVERTED_ENABLE_ICEGATE_PORTA;
	defparam PLL_inst.ENABLE_ICEGATE_PORTB = CONVERTED_ENABLE_ICEGATE_PORTB;
	defparam PLL_inst.TEST_MODE = CONVERTED_TEST_MODE;
	defparam PLL_inst.FREQUENCY_PIN_REFERENCECLK = FREQUENCY_PIN_REFERENCECLK;


endmodule
