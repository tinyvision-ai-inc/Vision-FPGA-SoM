`timescale 10ps/1ps
module QuadClkMux(I, O);
input I;
output O;

	assign O = I;


endmodule
