`timescale 10ps/1ps
module SRMux(I, O);
input I;
output O;

	assign O = I;


endmodule
