`timescale 10ps/1ps
module IpOutMux(I, O);
input I;
output O;

assign O = I;


endmodule
