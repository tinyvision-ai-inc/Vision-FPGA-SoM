`timescale 1ns/1ns
module AND2 (A, B, O);
input A, B;
output O;
   assign O = A & B ;

endmodule
