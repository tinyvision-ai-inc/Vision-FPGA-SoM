`timescale 10ps/1ps
module Span4Mux_s3_v(I, O);
input I;
output O;

	assign O = I;
	

endmodule
