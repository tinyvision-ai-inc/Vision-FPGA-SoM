`timescale 10ps/1ps
module DummyBuf(I, O);
input I;
output O;

	assign O = I;


endmodule
