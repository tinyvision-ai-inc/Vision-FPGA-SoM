`timescale 1ps/1ps
module VCC(Y);

    output Y;

supply1 Y ;

endmodule
