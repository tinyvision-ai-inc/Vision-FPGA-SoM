`timescale 1ps/1ps
module MIPI_TX_4LANE (
//Common Interface Pins
input 		PU,
input		LBEN,
input 	[1:0]	ROUTCAL,
input 		ENPDESER,
input       	PDCKG,

// DATA0 Interface pins
inout		DP0,
inout		DN0,
input 		D0OPMODE,
input 		D0DTXLPP,
input 		D0DTXLPN,
input  		D0TXLPEN,
output 		D0DRXLPP,
output  	D0DRXLPN,
input 		D0RXLPEN,
output 		D0DCDP,
output		D0DCDN,
input 		D0CDEN,
input  		D0TXHSPD,
input 		D0TXHSEN,
input    [7:0]  D0HSTXDATA,
input  		D0HSSEREN,
input 		D0RXHSEN,
input  		D0HSDESEREN,
output 	 [7:0]	D0HSRXDATA,
output 		D0HSBYTECLKD,
output 		D0SYNC,
output 		D0ERRSYNC,
output      	D0HSBYTECLKSNOSYNC,
// DATA1 Interface pins
inout		DP1,
inout		DN1,
input 		D1DTXLPP,
input 		D1DTXLPN,
input  		D1TXLPEN,
output 		D1DRXLPP,
output  	D1DRXLPN,
input 		D1RXLPEN,
output 		D1DCDP,
output		D1DCDN,
input 		D1CDEN,
input  		D1TXHSPD,
input 		D1TXHSEN, 
input    [7:0]  D1HSTXDATA,
input  		D1HSSEREN,
input 		D1RXHSEN,
input  		D1HSDESEREN,
output 	 [7:0]	D1HSRXDATA,
output 		D1SYNC,
output 		D1ERRSYNC,
output 		D1NOSYNC,
// DATA2 Interface pins
inout		DP2,
inout		DN2,
input 		D2DTXLPP,
input 		D2DTXLPN,
input  		D2TXLPEN,
output 		D2DRXLPP,
output  	D2DRXLPN,
input 		D2RXLPEN,
output 		D2DCDP,
output		D2DCDN,
input 		D2CDEN,
input  		D2TXHSPD,
input 		D2TXHSEN, 
input    [7:0] 	D2HSTXDATA,
input  		D2HSSEREN,
input 		D2RXHSEN,
input  		D2HSDESEREN,
output 	 [7:0]	D2HSRXDATA,
output 		D2SYNC,
output 		D2ERRSYNC,
output 		D2NOSYNC,
// DATA3 Interface pins
inout		DP3,
inout		DN3,
input 		D3DTXLPP,
input 		D3DTXLPN,
input  		D3TXLPEN,
output 		D3DRXLPP,
output  	D3DRXLPN,
input 		D3RXLPEN,
output 		D3DCDP,
output		D3DCDN,
input 		D3CDEN,
input  		D3TXHSPD,
input 		D3TXHSEN, 
input    [7:0] 	D3HSTXDATA,
input  		D3HSSEREN,
input 		D3RXHSEN,
input  		D3HSDESEREN,
output 	 [7:0]	D3HSRXDATA,
output 		D3SYNC,
output 		D3ERRSYNC,
output 		D3NOSYNC,
// CLOCK Interface pins
inout		CKP,
inout		CKN,
input 		CLKDTXLPP,
input 		CLKDTXLPN,
input  		CLKTXLPEN,
output  	CLKDRXLPP,
output  	CLKDRXLPN,
input  		CLKRXLPEN,
input  		CLKTXHSPD,
input 		CLKTXHSEN,
input       	CLKTXHSGATE,
input  		CLKRXHSEN,
output      	CLKHSBYTE,
// Universal MIPI PLL Interface pins
input 		PLLPU,
input 		PLLREF,
output 		PLLLOCK,
//Universal MIPI PLL Serial Configuration Register Interface pins
input 		PLLCFGSRDI,
input 		PLLCFGSRRESET,
input 		PLLCFGSRCLK,
output 		PLLCFGSRDO
);
//parameter PLLCFG_DEFAULT = 20'h00000;
parameter DIVR = 5'b11111;   //Ref Clk divider
parameter DIVF = 8'b11110000; // Feedback divider
parameter DIVQ = 2'b00;       // VCO divider
parameter TEST_MODE = 1'b0;
parameter TEST_BITS = 4'b1001;

wire BITCLK_int; 

X1082T001 u_mipi_txrx_analog(
	// Power and Grd Pins 
	.VDDA(1'b1),
	.VSSA(1'b0),
	.VDD(1'b1),
	.VSS(1'b0),
	.DVSS(1'b0),
	//Common Interface Pins
	.BITCLK(BITCLK_int) ,
	.PD(~PU),
	.LB_EN(LBEN),
	.ROUT_CAL(ROUTCAL),
	.ENP_DESER(ENPDESER),
	.PDCKG(PDCKG),
	// DATA0 Interface pins
	.DP0(DP0),
	.DN0(DN0),
	.D0_OPMODE(D0OPMODE), 		// Input from digital to indicate mode of operation TX or RX
	.D0_DTXLPP(D0DTXLPP),
	.D0_DTXLPN(D0DTXLPN),
	.D0_TXLPEN(D0TXLPEN),
	.D0_DRXLPP(D0DRXLPP),
	.D0_DRXLPN(D0DRXLPN),
	.D0_RXLPEN(D0RXLPEN),
	.D0_DCDP(D0DCDP),
	.D0_DCDN(D0DCDN),
	.D0_CDEN(D0CDEN),
	.D0_TXHSPD(D0TXHSPD),
	.D0_TXHSEN(D0TXHSEN),
	.D0_HSTX_DATA(D0HSTXDATA),
	.D0_HS_SER_EN(D0HSSEREN),
	.D0_RXHSEN(D0RXHSEN),
	.D0_HS_DESER_EN(D0HSDESEREN),
	.D0_HSRX_DATA(D0HSRXDATA),
	.D0_HS_BYTE_CLKD(D0HSBYTECLKD), // Byteclk output from Lane0 deserializer
	.D0_SYNC(D0SYNC),
	.D0_ERRSYNC(D0ERRSYNC),
	.D0_HS_BYTE_CLKS_NOSYNC(D0HSBYTECLKSNOSYNC), // This output will be D0_NOSYNC or D0_HS_BYTE_CLKS based on D0_OPMODE
	// DATA1 Interface pins
	.DP1(DP1),
	.DN1(DN1),
	.D1_DTXLPP(D1DTXLPP),
	.D1_DTXLPN(D1DTXLPN),
	.D1_TXLPEN(D1TXLPEN),
	.D1_DRXLPP(D1DRXLPP),
	.D1_DRXLPN(D1DRXLPN),
	.D1_RXLPEN(D1RXLPEN),
	.D1_DCDP(D1DCDP),
	.D1_DCDN(D1DCDN),
	.D1_CDEN(D1CDEN),
	.D1_TXHSPD(D1TXHSPD),
	.D1_TXHSEN(D1TXHSEN),
	.D1_HSTX_DATA(D1HSTXDATA),
	.D1_HS_SER_EN(D1HSSEREN),
	.D1_RXHSEN(D1RXHSEN),
	.D1_HS_DESER_EN(D1HSDESEREN),
	.D1_HSRX_DATA(D1HSRXDATA),
	.D1_SYNC(D1SYNC),
	.D1_ERRSYNC(D1ERRSYNC),
	.D1_NOSYNC(D1NOSYNC),
	// DATA2 Interface pins
	.DP2(DP2),
	.DN2(DN2),
	.D2_DTXLPP(D2DTXLPP),
	.D2_DTXLPN(D2DTXLPN),
	.D2_TXLPEN(D2TXLPEN),
	.D2_DRXLPP(D2DRXLPP),
	.D2_DRXLPN(D2DRXLPN),
	.D2_RXLPEN(D2RXLPEN),
	.D2_DCDP(D2DCDP),
	.D2_DCDN(D2DCDN),
	.D2_CDEN(D2CDEN),
	.D2_TXHSPD(D2TXHSPD),
	.D2_TXHSEN(D2TXHSEN),
	.D2_HSTX_DATA(D2HSTXDATA),
	.D2_HS_SER_EN(D2HSSEREN),
	.D2_RXHSEN(D2RXHSEN),
	.D2_HS_DESER_EN(D2HSDESEREN),
	.D2_HSRX_DATA(D2HSRXDATA),
	.D2_SYNC(D2SYNC),
	.D2_ERRSYNC(D2ERRSYNC),
	.D2_NOSYNC(D2NOSYNC),
	// DATA3 Interface pins
	.DP3(DP3),
	.DN3(DN3),
	.D3_DTXLPP(D3DTXLPP),
	.D3_DTXLPN(D3DTXLPN),
	.D3_TXLPEN(D3TXLPEN),
	.D3_DRXLPP(D3DRXLPP),
	.D3_DRXLPN(D3DRXLPN),
	.D3_RXLPEN(D3RXLPEN),
	.D3_DCDP(D3DCDP),
	.D3_DCDN(D3DCDN),
	.D3_CDEN(D3CDEN),
	.D3_TXHSPD(D3TXHSPD),
	.D3_TXHSEN(D3TXHSEN),
	.D3_HSTX_DATA(D3HSTXDATA),
	.D3_HS_SER_EN(D3HSSEREN),
	.D3_RXHSEN(D3RXHSEN),
	.D3_HS_DESER_EN(D3HSDESEREN),
	.D3_HSRX_DATA(D3HSRXDATA),
	.D3_SYNC(D3SYNC),
	.D3_ERRSYNC(D3ERRSYNC),
	.D3_NOSYNC(D3NOSYNC),
	// CLOCK Interface pins
	.CKP(CKP),
	.CKN(CKN),
	.CLK_DTXLPP(CLKDTXLPP),
	.CLK_DTXLPN(CLKDTXLPN),
	.CLK_TXLPEN(CLKTXLPEN),
	.CLK_DRXLPP(CLKDRXLPP),
	.CLK_DRXLPN(CLKDRXLPN),
	.CLK_RXLPEN(CLKRXLPEN),
	.CLK_TXHSPD(CLKTXHSPD),
	.CLK_TXHSEN(CLKTXHSEN),
	.CLK_TXHSGATE(CLKTXHSGATE),
	.CLK_RXHSEN(CLKRXHSEN),
	.CLK_HS_BYTE(CLKHSBYTE)
);

X109T001 u_mipi_txpll_analog (
	.VDDA(1'b1),
	.VSSA(1'b0),
	.VDD(1'b1),
	.VSS(1'b0),
	.PD(~PLLPU), 
	.TST(4'b0),       
	.CN(DIVR),
	.CM(DIVF),
	.CO(DIVQ),
	.CLKREF(PLLREF),
	.OUTP(BITCLK_int),
	.OUTN(),
	.LOCK(PLLLOCK)	
 );





endmodule //MIPI_TX_4LANE
