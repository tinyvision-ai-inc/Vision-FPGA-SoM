`timescale 1ns/1ns
module I2C_B (SBCLKI, SBRWI, SBSTBI, SBADRI7, SBADRI6, SBADRI5, SBADRI4, SBADRI3, SBADRI2, SBADRI1, SBADRI0, SBDATI7, SBDATI6, SBDATI5, SBDATI4, SBDATI3, SBDATI2, SBDATI1, SBDATI0, SCLI, SDAI, SBDATO7, SBDATO6, SBDATO5, SBDATO4, SBDATO3, SBDATO2, SBDATO1, SBDATO0, SBACKO, I2CIRQ, I2CWKUP, SCLO, SCLOE, SDAO, SDAOE);

	//Port Type List [Expanded Bus/Bit]
	input SBCLKI;
	input SBRWI;
	input SBSTBI;
	input SBADRI7;
	input SBADRI6;
	input SBADRI5;
	input SBADRI4;
	input SBADRI3;
	input SBADRI2;
	input SBADRI1;
	input SBADRI0;
	input SBDATI7;
	input SBDATI6;
	input SBDATI5;
	input SBDATI4;
	input SBDATI3;
	input SBDATI2;
	input SBDATI1;
	input SBDATI0;
	input SCLI;
	input SDAI;
	output SBDATO7;
	output SBDATO6;
	output SBDATO5;
	output SBDATO4;
	output SBDATO3;
	output SBDATO2;
	output SBDATO1;
	output SBDATO0;
	output SBACKO;
	output I2CIRQ;
	output I2CWKUP;
	output SCLO;
	output SCLOE;
	output SDAO;
	output SDAOE;


	//IP Ports Tied Off for Simulation
	//Attribute List
	parameter I2C_SLAVE_INIT_ADDR = "0b1111100001";
	parameter BUS_ADDR74 = "0b0001";
	parameter I2C_CLK_DIVIDER = "0";
	parameter SDA_INPUT_DELAYED = "0";
	parameter SDA_OUTPUT_DELAYED = "0";
	parameter FREQUENCY_PIN_SBCLKI = "NONE";
	`include "convertDeviceString.v"
	//Converted Attribute List [For Device Binary / Hex String]
	localparam CONVERTED_I2C_SLAVE_INIT_ADDR = convertDeviceString(I2C_SLAVE_INIT_ADDR);
	localparam CONVERTED_BUS_ADDR74 = convertDeviceString(BUS_ADDR74);
	localparam CONVERTED_I2C_CLK_DIVIDER = convertDeviceString(I2C_CLK_DIVIDER);
	localparam CONVERTED_SDA_INPUT_DELAYED = convertDeviceString(SDA_INPUT_DELAYED);
	localparam CONVERTED_SDA_OUTPUT_DELAYED = convertDeviceString(SDA_OUTPUT_DELAYED);

	I2C I2C_inst(.SBCLKI(SBCLKI), .SBRWI(SBRWI), .SBSTBI(SBSTBI), .SBADRI7(SBADRI7), .SBADRI6(SBADRI6), .SBADRI5(SBADRI5), .SBADRI4(SBADRI4), .SBADRI3(SBADRI3), .SBADRI2(SBADRI2), .SBADRI1(SBADRI1), .SBADRI0(SBADRI0), .SBDATI7(SBDATI7), .SBDATI6(SBDATI6), .SBDATI5(SBDATI5), .SBDATI4(SBDATI4), .SBDATI3(SBDATI3), .SBDATI2(SBDATI2), .SBDATI1(SBDATI1), .SBDATI0(SBDATI0), .SCLI(SCLI), .SDAI(SDAI), .SBDATO7(SBDATO7), .SBDATO6(SBDATO6), .SBDATO5(SBDATO5), .SBDATO4(SBDATO4), .SBDATO3(SBDATO3), .SBDATO2(SBDATO2), .SBDATO1(SBDATO1), .SBDATO0(SBDATO0), .SBACKO(SBACKO), .I2CIRQ(I2CIRQ), .I2CWKUP(I2CWKUP), .SCLO(SCLO), .SCLOE(SCLOE), .SDAO(SDAO), .SDAOE(SDAOE));
	defparam I2C_inst.I2C_SLAVE_INIT_ADDR = CONVERTED_I2C_SLAVE_INIT_ADDR[9:0];
	defparam I2C_inst.BUS_ADDR74 = CONVERTED_BUS_ADDR74[3:0];
	defparam I2C_inst.I2C_CLK_DIVIDER = CONVERTED_I2C_CLK_DIVIDER;
	defparam I2C_inst.SDA_INPUT_DELAYED = CONVERTED_SDA_INPUT_DELAYED;
	defparam I2C_inst.SDA_OUTPUT_DELAYED = CONVERTED_SDA_OUTPUT_DELAYED;
	defparam I2C_inst.FREQUENCY_PIN_SBCLKI = FREQUENCY_PIN_SBCLKI;


endmodule
