`timescale 10ps/1ps
module Sp12to4(I, O);
input I;
output O;

	assign O = I;
	

endmodule
