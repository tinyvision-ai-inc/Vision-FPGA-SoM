`timescale 10ps/1ps
module IoInMux(I, O);
input I;
output O;

	assign O = I;


endmodule
