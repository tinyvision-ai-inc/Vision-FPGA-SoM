`timescale 10ps/1ps
module Span12Mux_s9_h(I, O);
input I;
output O;

	assign O = I;
	

endmodule
