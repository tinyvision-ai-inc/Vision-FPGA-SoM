`timescale 1ns / 10ps 
module SVSS_sbt_a ( VDDIO );
input  VDDIO;

endmodule
