`timescale 10ps/1ps
module Span4Mux_s0_h(I, O);
input I;
output O;

	assign O = I;
	

endmodule
