`timescale 10ps/1ps
module FILTER_50NS ( 
			FILTERIN,	
			FILTEROUT 
			); 

input FILTERIN; 
output FILTEROUT; 


assign FILTEROUT=FILTERIN; 



endmodule
