`timescale 10ps/1ps
module PRE_IO_GBUF (	
	GLOBALBUFFEROUTPUT,
	PADSIGNALTOGLOBALBUFFER
	);

input PADSIGNALTOGLOBALBUFFER;			
output GLOBALBUFFEROUTPUT;	

assign GLOBALBUFFEROUTPUT = PADSIGNALTOGLOBALBUFFER;


endmodule  //PRE_IO_GBUF 
