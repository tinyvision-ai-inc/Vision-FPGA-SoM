`timescale 1ns/1ns
//The following SB_* Special Primitives are broken due to many of them having
//integer parameters assigned to underlying string paramters. These SB_*
//primitives are needed by LSE for legacy code however, and LSE will take care
//of the conversion from integer parameters to string parameters.
module SB_DFFER (Q, C, E, D, R);
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Lattice Semiconductor Corporation"
`pragma protect author_info="Lattice Semiconductor Corporation"
`pragma protect encrypt_agent="Radiant encrypt_hdl"
`pragma protect encrypt_agent_info="Radiant encrypt_hdl Version 1.0"

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP15_1"
`pragma protect key_method="rsa"
`pragma protect key_block
ZnOtAiM31nxJOxNI2cd7Lt85oD8uBT0RbbbYPfQ/Q4DwlP+61gLH+wrHpiCGQJaW
Z8teUJ1JSkcbccvl33JMpTxuxHWyuOplDch4wimltRfqxz/wwfvxzEKHKTq6iA1s
GwZ6Codnj11D+vQUffBVciFlXYOH3U3S3br9oHEDhfC6Ak593KKowcfOYV6dFs8o
wAt91EYOCwejJjTX37zJo21B8JumEV5NBZJOHlzoKvAJ+txESVViBtgP95pguzEm
1Pq2Ys+XCwronw6zmLREJVA+Kdu4hIH00d11xwine3iSf4ALNO6M+Gkwy0DyaULp
OF+yCzI3jLTDVPX91hdvJw==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
LPpc4I4yQFHvIofyx0vaRrAA8DQUfZG4xLL/28HZ3dIwrTMZQtWgeGIenEmigE6J
3Mo3Msba00YsWrmJmCmnTAT1keDk8Ru9Y6N3gjPNH4M6EGKhLNmNPQ7D4dcU1ZuC
YqVioNAc+m+fTosOiOlqeOxhUfaEfemWPJ5S6HhXcfJEyegAhfHFfnhpoPvDsX3+
NzVoIQePFbFNrJMRAN/PaQwhnIBchb/Bby94faTWnj4skjjfMXB6QtY1jM7fBngk
tW0iESGtXVwJGMnXtbm6m060EylIh1fRB6U83djn9gGEJnbezWz2lkTAGQMB236p
SeqbomMuRjSDzdH/qxUWIQ==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-2"
`pragma protect key_method="rsa"
`pragma protect key_block
qkJaZ9XHw25O00tXnY9NgBF197y9ZwVOd6xAAuKsKpNCYcQVwrxdAkB5Dxq6YMi+
M2Y1we+5S/vXoZGvNhxyn3uNJ37zhdKTgH+xd0jwkn6IzAp4oiICaRfknmne68vO
40I6eLt5zNuQWGKK2LiRgJZ9+7UcsmDwSdop7C7syaNxkBgVa5irNEGvDdexucM9
cFmW/17ufJflZvqQ3sRw3Zg33xjWVAlTIxitarSEUMx4kR3RIvo3RnTAHQcfeJAP
4KzG2CKxhZ4Ro4PXjh+t8ZvglM+nwRqJNERWvxXSq7jbE+5uop8g/PlSpXBhAF17
x75Zfi29v2nVUL/AzlBD/A==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=128)
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect key_block
LDQi+MsfcqLOBDetUvX1uKDt3Rd+JEEoCYh8yDhtHqtjkFyMaiZ7uJbdW5461JW5
INnz7hn37E0jv7I4LQX5SMNT/96NrSBOg47nu0vAc5R097eMv5EG+Bfbs2EYQzPG
6koi/IP9lJs//f28lfjmvy1uV0NRQU46NNzGtblmWbs=

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Aldec"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect key_method="rsa"
`pragma protect key_block
vrLhfBc84ZxhpOVDydPCueYr8R053VUGKMGbjqzyqtj5bhA8oVSQ0uB/J4H7OA0D
Ou1U6/HmICZAezP2ZlwKnkz75jh05EPXbgRIvOWA4ljL3wjOyPZfpVdg5Wca3LYj
2Ep2GZN5mUlKpMiJpCpu1iirnHB6Axw5h9l9CSe1pWnUCQhMSnx3nYMcgSqcbnFZ
1BJjfmiaGZtjmCpwOU2lwyEkjb0jfCryJ1pXKXNf6x5qZ1p3l7Pt5hde70aUh4Mf
oHWsjo9x36jfdmfdcROR4a/Wj1Tctf0pgTfMY/M96JeKSjHVUHVAM5010PqY9/Zy
vgLcIQ2VRxw6+vpUXLGUvg==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect key_method="rsa"
`pragma protect key_block
pLYSqQSsSNOeeDWc956mJQAm8AikOQE2GcnUdQ5KdMh4RbmdAXQkXOvHT+1/PXyF
4+3bw3UwDf8WvEG6UOLMfybQWBVfOHzu54GuX4/6l4ct6nFaLQQdKlCs5T10DPm7
lIrIsKFwNT3DdZHE6VEUvDFdoJvQQydbrBNlxi6hMdj6rKA3gy+whoHFNxFOsy1H
8EU6njLZ16Mlu02UKUZPwUGmb6uD9owQ352hoY9mBv/HZV4Xft1LLKNXPXg5VdWY
2CgNm5qIBMS00Li+0u3s7t3yP0vq/tA+XHrsujgP0n8ivmHciOsnqcVU7D49PMHp
iisqpEabPqJvut+lAX2NcQ==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Lattice Semiconductor"
`pragma protect key_keyname="LSCC_RADIANT_1"
`pragma protect key_method="rsa"
`pragma protect key_block
lzgFGcgFAOpaGWSEXLkjKjbOp9qBt7PYXrWI+woAUxL0BooR4pS3axxtnuHoL0oR
/XqFKV/p4kbO6nee9VUFnFgB8W4zIELoUqwhpeIJP2Qye1GLPjURopikq2qZNrb3
kV5+sSxApHBFdn+Tsy8TM5Y5CNZM4X2VMh7d658gW3mIFUn457wBOgfx8U+T9y64
AoQJFk8wNnHeeLhiIr99yFh9rJjS/jSWGbdsDdDrvmbOsvwCpkE1I72E0lA12b84
r8bJFgsfAVrGeC6oHrdFbXm6ogZTNI4eSSpT/JPwg9kQFUr9FtkwznHusf2atM7F
LCmEoxGnO0/9/jS4sKIQ5A==

`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype="base64", line_length=64, bytes=176)
`pragma protect data_block
thtmAmZ9zjuCYUmc70LI8x0788xtKQPPCvBY4anJtHPAAPochqIMg6M99f43zvDl
O9amDRsm9vrl43yWJAIeNxNlZKGlBL6+5HoFWFRcubyScXpTGr+hkFLvKc3U4Kr2
ocL/5TUWeXYVQy9b65vm7xCSapBl7aP8u0T/haOKm5fkyiPovttZu+7viCtDY2Vc
ZxKqawDUUct9T9ticq6XT1kaSp13c1rTQaicSGDjMaE=

`pragma protect end_protected
endmodule



module SB_DFFESR (Q, C, E, D, R);
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Lattice Semiconductor Corporation"
`pragma protect author_info="Lattice Semiconductor Corporation"
`pragma protect encrypt_agent="Radiant encrypt_hdl"
`pragma protect encrypt_agent_info="Radiant encrypt_hdl Version 1.0"

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP15_1"
`pragma protect key_method="rsa"
`pragma protect key_block
iPL20x68pU/oVWhRt4QCqbcVYdX9iU23qbzw0qFqzn/fyaS1jV8iTI717DesWN/m
djX3bQUKE5smdFSlNTysRpNDq4as/vGKTSdVuM9y8Pv+qr8OPrZeTOKVEEEt1JKA
CiUE3uYT8ZYM/lUgaBdCVXJd8J3LtC+G9TzTSOhdWEew0a5BgXztO+x7FSqCvSNa
7E4h7qdGX5tPOy0qMAFJwHW8Z11kpA2x5XrT4yLwQB8oKo81hlP3aOAHLsJM50lV
Gdq3qHdWRo/vXAoMxQlC3j7reuVDZBeKE5n785z4w1Yxmr8zN5TMZxeYQH8/9y64
ppSsx9k0Tiinky+Fh0V9bA==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
rVEuGd7JSzf62kQiVs7SH2A69swfJe8grCqHtLDT8sGNN51+XZrniYB8g4idSL2w
d75bcJPN7leJ6flcbvN7Ur/1iTihuORpJ7owYVSuO9NIv8OSnOtW9/QgbziCJ20H
JpX+KBfFDxv5cYvhAcYIcOFaldNPUT4AvUS/MfiN8Pvyf4BQvz2lJBQtPraT5vgM
gMvhDX0McDZkerIenEYHWyW0qVyvRckrK34SI6rRWcuXgKEfK6ANU4Qgb6gd9K5r
VTOcNYXQ+WXgr9gnaBt0hFvVQRZtxC4J71JXFS/eEqCnfGrP2vRLIZxcZAyeubVM
L/GfTPfFtEgRy0RhK4iRVA==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-2"
`pragma protect key_method="rsa"
`pragma protect key_block
Xe/AW48ZMBwTyqYBx4j7Z0upFJikfH1Cj/FRk9rUzqDiO1a2aXlv9UdKegCdUPmX
OFNDeFU6qCAQ2IIeCnoqTDVCfeklX9L/XDJbDnrXPK3bmd+AHlYGsEkMfZpUPVKv
e9CUQF2lLym3eDzqmFGFMLdJlxYkCDRZHfO1caaSqxcC1pMo4+1ESAwm8QrRPAKC
ncILv0hiA9GwncsYanH9TgrHPdPTa7UCplQrvaEZQAks9c8hM1L3c6ouA7tZxHB3
SK7MTfD0xkfjakd6luN3YlbwQDes2WEKXkzzOrUV/L1PK9iXee89mb1BQTtPYHzk
SLd3IY9yF+X8YHLs8jk2Sw==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=128)
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect key_block
1LX+3DDXjtCMGeN3O0IQpzsLpOGa2fii5qRRplGCJz4lAd6a3eI2BVhbrj4Tw2rR
girl/inNY/BIyT5fT/P5RLQoZjZ4RbwyuNEBNdmAxFZzD6AUDtrTrK/v6D8pBjx4
EC61fyQ1hNR3FN4WXpQ/ytIp/5KppvvHV50lNxqRw30=

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Aldec"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect key_method="rsa"
`pragma protect key_block
vrJmRrdIetwpR9JGaSQq3w/KvsohzUktq4ttZjX0QYleU0KC3rccULkVyav6793C
NJXuMMcNzFEC5gQNtpJW9EtsWqiBdLdXqXylD5cqOWGzKzXQ+t0JztzC0SsOxGCS
waInJC4DlEEUiQCrai35STZmSeRmT+0jx71/4AuLxC53CAQBqkZQVWLPfs8RUq9j
NOxbOghyoD68xI0ys5TsOi2TWLl/TqeVe+opONiQHO/udFcXyeQcLJa9Ah8lJlYm
XjfoE4BfMZ9Nu7kUg1OFuJJM0TV9wqn8d+HFhbdXn8+aymvjACGcgypYbfCbtSyq
2sn0Cn3kgG3zfYUDVjAB5g==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect key_method="rsa"
`pragma protect key_block
KaqHyZdJedEsE/jw5q/kh/Rw8w0gLppZjLbdkI16H76xmSZyxsobIuTZvOkQJ357
U/lU5i2QsfR0YzqCd0LjrgavWp++EMy7L+sf0u8ZHQBmhgHkKA6glM4WnlJwMaLh
DoqVtv/iw3S26/iBzu2YnJGdqqID7yeshtWE6yiU5+IUkrpMD+vk2cwTWJbC/3Cm
fk5Brjgm37gyvqvJwbr83tXZV+7uURLy3QG2jzf1bLiurQocstXWCydiXMrzeLPw
155KZfKX2/bcx7+czxaQ1lFBWJ8+HyB6c7JbhgWnasVHVxLg91SJ7R+gA5f+dieX
JNMltzYMHGgZBU85Gdb+bg==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Lattice Semiconductor"
`pragma protect key_keyname="LSCC_RADIANT_1"
`pragma protect key_method="rsa"
`pragma protect key_block
fyCOz/yZt9ivlNDGZZ2KQp2PnXCtQZWC+TnikkpHl4AyCIQQKyPHo88UVoQSUyU+
uH737k9QBQyAsv3MUf9yZ3PgdEtqfA+kazt4Lv+P/TxzweL6rHCM6ay2geMgbvww
3BdFh0FOvYPMX88PO6+Zf1zp1E9QIuMbl8fgazQl4k72dQG3L4nSyMkL/XLWEit1
2rNOiZeloor8vGCYu+opJYi/7MbS+7IVcE2GrDm0k56mmKO5q4L7p5+HlcSLSaJD
QnpzHNn8a31hEBCsvh2LaRE0IrTzB2CCvOyRqDoUT6x6MEfHoIA0EblF4f5K16vc
HF6iirCNjyU73VsKbbGFUg==

`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype="base64", line_length=64, bytes=192)
`pragma protect data_block
hAV/ADXJCn+8/WUp+1eaEfnh+ghqiO3fV1SqgJYAX5nNSbSCrm+bYjtV/QmruqWk
Y+kdxddJx5zGb3j1yUIf98jVdcd2Qsd4qV1B+b5ftjfUCZ84I1BOeJjMMJL/BQDg
zmYpO1F4OFphMvj3GrMJRJYnN5XGklaWM+NPJOLcfijodGE04Dev/k0TxN5JK4Yy
J4Pm9VwI4KrafllzdHZF9msyr8mrgR8mQhNsX9SlWA48hppl/CYjtpFsV/RMEpzY

`pragma protect end_protected
endmodule



module SB_DFFESS (Q, C, E, D, S);
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Lattice Semiconductor Corporation"
`pragma protect author_info="Lattice Semiconductor Corporation"
`pragma protect encrypt_agent="Radiant encrypt_hdl"
`pragma protect encrypt_agent_info="Radiant encrypt_hdl Version 1.0"

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP15_1"
`pragma protect key_method="rsa"
`pragma protect key_block
6BbVRC0c25AeIh+E0bNjVoczsXqnJdQoYWfElziIRV0DSf1lA0ZgWV45xnEDXqv3
NhHQ6d5OGu4wjKjhdSpKf9sbiif53KHiez6k+ySn/DgbiZm67z1qK6SHWMlynyFM
guDP04Ym9P0XIQklgOmmwv87lrLEbwTqktD9fwBP0WHyf1kYT8Mm8EYCj4LRYq65
l8cdogcX0JcYktgQGGmZ47/SjHZoo/dkZy56Y2HRtQlBXcqlyTr5t/yBmYEU/qWv
IJy/AEsVsxTpqSw20UgLRcv2oxk/yOr6lZEvyzI6T3DwrtBSWf3xGawexWixWPi4
d67976wKTGcEDh2l+vghEg==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
GX4f9G2xa7q5lsX/mMmR0mX3rMW1KEUAwoKX3q4Jhmgz8KlmVaFer41YuUYsaKps
Ch1IKvvD2vif0ApogGFIyBA6lL1289lC/kiju8yNN8Cf771RGvKKqRGfHX6ayqJE
NOCYBBxfUjdvMFu5FZ0teFsM+dUh0zMNl2xheJXtZ8pdVRO0wLDkbTzHVOyVte+7
jr5QHI8Ii7m9TrqxV07OvmjPuoxVUxueiyNk5imO2w2hlwrZVSX5bzPQQpm0sDps
jUk84Ie+y3J9rzUFpOE0asD5xsZu2CBmQwvxczT4gWs5CNzzvVlDcVgEAAUXr1BD
oHdGfDy0aKHojTq2JqEtvw==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-2"
`pragma protect key_method="rsa"
`pragma protect key_block
LjIb7F+z+7UZc21rLjqL8CQLEdQFf22zZbASobKCIkglSwxyU7kcqtq3jBZ2HLEI
KWvotWeJTnZnIUPBYy5YUSNotfR1Vh1L+PKSfouqyNLmYDxL0N7K2ycWMQdokXkN
qKNsPJbrIEWVlVedkAT8UoLvP43oE+z70l2WOCce0ng5xAhscAZMWiiTz163S5R2
+2nyU0u+349439ZwDstplZA5fTAULNxxpPzXerNHW9sVjFqVRKrLhoEzeUSFTwRG
2zUfAEg0DOY6yWrX60hv7bFpROpiLn7nyWgUFNQgYghvRdhqVQCvfDotFNg8EYrM
DWIy9acXbPzXVPzVgrPS7A==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=128)
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect key_block
Xy1chi8geKCeaK3I9x+MfP0y+iqorB5dL5wYdpn8AKzayQ7ZceN+q49Zw6zprcZL
ETznerJEBzLcjrA26JBFfbYdJ8YAvmAaa4nVg+Ql3QMizQcscMH2gA8RFqOiZv82
sy0fXSp3HSvx5ye+gmzfh6ZcZoX+Y6nuQ3npRZw84VA=

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Aldec"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect key_method="rsa"
`pragma protect key_block
miGWQfjXwXcNLjTySsFffC98mJmrrJn3+RBlqJP6hJP6XqaJDMl2bdNcghzLj/kt
SDFeEafVXQa9UCM9PvCasQZv9/3TDkuTlwsflm2Ng6m8VgDWWkqz/ag9STu/IAxN
AefzFjgT/gzyVFNVbm3T+ifSGnmxCkFg+Ux9XXPvOvj0jgNPWPgMHxD+elhHQAMf
k2FwdAkAQya2oIp/JbsxT8nY8BSXxXeritoHIVbEnf00SP+xF5nEhDGw1VBkbUYY
ZpVG8WlLAw/p+o3FzinIX0ncUEfDNOInWzf9ChGJL6BUP+rpbEIfe50SYKROu7cd
FtkEYbd+Ru/oJ97StMlGQQ==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect key_method="rsa"
`pragma protect key_block
jLDcphiYovtsFU9n+aia3BWOAiWU+AmCYA1OuLXnjDGcNRyJcsB2OywZh9C/VYxz
qCwqlmku4JayyOJpFwUAftv4LLdmsfYkkw1hdJNngXY64XMh53E/Acu4b4qFHx1N
JeZ34TCdV09D6miT1suC2Ux7xAcErJ7RuwCnCsGCC5dnPQNQAoEqgMR5Y/53rVJH
9MGVAtroPGbm3qbaiR4WwU7D3f8igUl4w5LEOc9GvsuiM3Paxb9qTL/Qe0ml3LGv
8j/Fn/Lqn0wAuSnm+3JvreqxZo4n6CgsE4kAux1FdhMWs0m7phcp130v45+mvqG1
OPX8HJpEoqyiJ14WYjPT0w==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Lattice Semiconductor"
`pragma protect key_keyname="LSCC_RADIANT_1"
`pragma protect key_method="rsa"
`pragma protect key_block
X9JTNMaUOJoDi1I3sNUXNxsWzybVCa2A5Oicnc4GnwYifgEedQspxY/CzQL3j01t
+JTds3s17RsyTV/ESTjp3QmNAzXhOF5cdXrylwvlCMRFu3Kg+epaeGcj8z6GamaM
ZZiAXB7+Tw2L0lmgT+2o10bh8twAoysCbXNC4jufTXLMAKlUIb3+QKweFzoTl/NN
LCsamOzcKefg9qA7sxT6bGFyqKXxbWz/XUd9+RJpVE2GQdhS6xvCWKs80ciwu8Sz
QLizacopixA9t8kYZZvUWwF3nJ8+h6eV6VKWNAvOFKWpa1o9y25MU0Q3Yl3r37TS
fzKETqVgBIDHOAzTCbpcew==

`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype="base64", line_length=64, bytes=176)
`pragma protect data_block
yuR7dda1FTUMMH/hs0U8H4c9qJtp/R0+3uRVb3inoBYNbdpzyRcd1wZsjyYuknmd
zyhn+3fUMdexzA3sc29LYQhxh87/9ydg9fbDwN6072RSUnv8VndwhPEXJ3NHrCJL
FE8RXhi9Ri9C4gS/G0jwfU39GXTid9v5vHEgnHfRAteWvKFDsSWvxvu3IH0tq2Qu
U+McZu9qG4ccfkM9GSjacKbVT8BAZvujWVYfnVKzyK8=

`pragma protect end_protected
endmodule



module SB_DFFES (Q, C, E, D, S);
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Lattice Semiconductor Corporation"
`pragma protect author_info="Lattice Semiconductor Corporation"
`pragma protect encrypt_agent="Radiant encrypt_hdl"
`pragma protect encrypt_agent_info="Radiant encrypt_hdl Version 1.0"

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP15_1"
`pragma protect key_method="rsa"
`pragma protect key_block
t77Mpoczsx6yPAnb6Ndgv18UO68WYsXZGFPEx0iJeIZNvq4RHDxdGNMSTTbdd57L
t+/mjRM0U2Y8kmOglexw60jhZdOppwub4D2U7Ucp3QaHVG6sAh/k5o4948qGf40D
SNCDu+wHWwVBKD6mTsei1rh7NHFOaWjiEVZkmBofaD4qe/cI3PUcmPE0dwtkA0Gw
6+tab6tnIh6lAmEiiYH/9EoXLvHzPp1r1lgw5LdETpUjGDRsdZStn8OsV5TuTX4u
53p+QbesgrnwnF5ySCp4HACte8bWPqUMVAxytwyaIOynqITc01Y6Coo+pkmD0zP3
mZ/4P9kWvgyxPjsoD2o3+w==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
QhvNqTgcSVlP/IGjpDtribuPu+KHLfp/kfAdblDRAEAyrILiBgrpNKGFoWCUSPjp
e3a4UcfqpR1xaI5ZrpyRUUZMN4ixgg7oLa7Gb7kdPWW+kuJdcA5VxrbU1ohHcJeI
+7oq4VbK1UcG73RYXGFJOYAkH0Bebx6kplbf+LzvmMLaprqQjcw/wofg2XrChPqs
D/Zzt9rX4YyaKmfKWeEJjbqLbXNCnMuTc7OBV12oipK6wv0zyM+JcL8lvcY1qBUH
Oodf8qlweA+5DZm6+79j94arBslbLNsj18E91zJHYUQdxRmlMLGcywJNlt0G6whj
+SK7e5q4uVzyPGY1bQBIpw==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-2"
`pragma protect key_method="rsa"
`pragma protect key_block
dSp9unAQQ5tNXv3YYvM/mfuzLEp9uW0aaM4v9mnNIUNESFUmlEnT0bg0FzMnz48m
9CjywTEI+fgu5xMAnyat/YIELL2Xf3natNf0QJphBRujM9S1WFNWCH4xKygWAf+G
v+3TiwsGUZ3Ycla5lV2zQr9yeUCP80HLSKrK4mmnbbkwnWLMxQreIXToW7ygIIAn
lvCd6oBqOFExK3sJTSrcHo1WsIEokjlPNEgfBpKvzKIqNafrw6T61vnityuhre1d
RbDs1BadkpZjzI7++3wf9mU1FGcf5mOEY5ogn6NTBjfBqfMYuEn8s6oITicoVnpf
O4P6g8xgnchk5kc8Ji8rWA==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=128)
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect key_block
AX/cdITaPuyvw7dCNDZHylY1GAqPUQNAe/IPqjVLs1Jj5rBSp+/VF/Sked/Oq8jn
6opAB8EPfe5euf56c2Vz9yJEoPYej3wHeVIa5RWPUI7zgKqVAipp5LvcNqRzS/gg
LPbA2exHsFd+Fk1fg9NMUt9u1KsI01KH1lxRq4dTDcI=

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Aldec"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect key_method="rsa"
`pragma protect key_block
LIuCle/zrl8yu17kRWxu3Kg9ayLeQTotGy4Z0ejjyt0Q+gXz1kAHpHy9G67smUR7
U7bu5S5kiTOA+uny3DZK/FWoJLzJb1AtC7XPg9GsShxnUtSCr9aONPD8FW3YZUHe
L+gTtl3kUWFbQIGBwh1FMBUhKEskodaqyIkVuu8RCRCs1D+ZoWc94VYfXoDhmzVv
rk1GCkvZNRahR8hKMHHEuX7LZYZgWcn5/JB4uzzKiDjM+jx4UblKiIrpe62IEwfI
bN0n/ckUHAkJ7dAno/yGr7g6lLM0lJXtuKOIywCqJc+xFfaIzIng1u51sLy7ZD7T
fvbNRB7ifQ0y86dTk65Rkw==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect key_method="rsa"
`pragma protect key_block
LQv6rdgxFvc/4/tCYRnNIqYEgLKrRCZQufYIbtHiqDqu+xn8cOyB/YNtB1x2J4pU
zLd7OKFnd+6fMZRBTQ4+1u223axCCD4Hhsi8e410qyat8zzoSFEtKi26dLbU+oDw
ItVOIb5PtGGODcA8DC34l0OkJgMlF8hlrKAhPJ3xV5cYW/IeBe4WhECKsY+tLI56
IVHwGGNpY0VoaO/t8ZBf4sC37M//bHN7FM72lh1AnIKlzOVS0HZ6XFDOeAlyxBeU
yHHCr1qACGVBZtbzyLqjjBTnCk9thIAWsc0gL0mX/CNDKi0F15mjzl1Z1C6pREAZ
qqtg6xIA5MZ/hTZxEuD4pA==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Lattice Semiconductor"
`pragma protect key_keyname="LSCC_RADIANT_1"
`pragma protect key_method="rsa"
`pragma protect key_block
CnM+qwKjnIfaV6JNiyl42ExZO+RQZBJGGsmuDfj+0BqyaYfvzYe9g4tasJeCm814
JJn+DMdHuU1ylLQz5B/1wYcgziLEgOqwdYRs8nJhzSOz+hr7+AGFteZUlrGrxlBV
PeuaRspO8mYFuEfUl5JpVGz0mT6R3JUvCFOh48r77YAmWfHCWGybuthTDMz2O6bS
3IKx5EmgZx06zueOLMOee2yn2pIpKn+IFKkvKQNXdteSYiESLxlE0PIm6eBR55S/
0MQ3hPt/zPN5EPgSr+lnFdjVOBNtDk5ZPA1MTSa26pMU5Wilk2rKbDvxigdT6JNo
+VH6p8nZ5vKXRTD/YtZW4Q==

`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype="base64", line_length=64, bytes=176)
`pragma protect data_block
T7lvXKXTnSl4QLozQ1N2TXshnE8WsIXSBXSfSifbc4aSeH+UDACFS7oBGZ8dnvEl
EtdaSPSrDUbUntQghOGybFCp8mpRXsBUhOzEgTa5BsrunYOcKd01vRHSiY278Z9y
odN78MXqvLFt7Yu4zxpR7H0vE1vmH2o9lhBlwU6UQabqgdipjMiuNJga00SO4z07
lG2O0mIdmb3kNvXzDVTkttpji4jQSqlzQ6tR91Oo+lM=

`pragma protect end_protected
endmodule



module SB_DFFE (Q, C, E, D);
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Lattice Semiconductor Corporation"
`pragma protect author_info="Lattice Semiconductor Corporation"
`pragma protect encrypt_agent="Radiant encrypt_hdl"
`pragma protect encrypt_agent_info="Radiant encrypt_hdl Version 1.0"

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP15_1"
`pragma protect key_method="rsa"
`pragma protect key_block
HyzfE7JHj08FY+ylkWdFQ7k3EiWwYjDU/ugeVtv/SAjID8FvkHjmurfPQl2zpTJA
k6EoaWUHVsWjp47nAVcKOaAObnAN+f450rL+btuk9tKayt69kXNwC9tFmIIgkHZj
Ww/wr9dH0Ib1EKIXAw3c6ieiJ95TaUuMS97d2vdVR0daH3HffV998BvWUUEXVQJH
oudQrbKOV32ES2qkmJbKGfnSlLwyRalkx5V8NhwHoaF3YfhjkIOLq5F27Zk7Vmrh
+DVThK/qZmk06yairK5jI7+QHIWTzUkgmfOrTUFn2o/vLCzUdM0q3h3IVED4E80u
c6Fwx03hZbViilxt/MrR1g==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
el3vbcT2c2RRyBL3+T0eqMHqz7G6yfYaK6l2wd+PDRWKs6VZfdw3+O1mYuDJuSvw
FpxEHC0z62oh/KdwEO++iuVy5Ie7mttzbUpziLkzE8/zS3uxZlbSD+ovUImtga1d
yyug7ayYTID8/MJR74hXQLGPio1Ck5LE9+O5Y+TCc54LnKYnF2IIr4MMTWviWemb
qzKg4y+qAIpSleUedx7eoGHcO8UMabFprwHLXnK6qvkSwWgQFJ2H8OAaFsAyUojQ
g4rId62/lsea8SU/Omj0WSm5verjPPZRkyT1zhFveeFo+7S2DzZfunZhcES+ecoD
Ahmw7XKjDNGz3kj6kckoxQ==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-2"
`pragma protect key_method="rsa"
`pragma protect key_block
oCZy9SZMm62OwhV5KaOMv3HVukF6udkrp6R5Kh6t4kaxz559WYevmrqW76ywUthm
Os3ZPq7ihDyD/pglRQhNAYKdihuHqjUykFzmvs2wD6PC1CVR7J71Ya/uiW/oS7RO
drq4XA1era17SLJO9Sn+pgTQhmhTJMSKMmUok28bjnitswt4xlCn++d1AGWDyV6T
3utIi42LFfXRHRyaLNxIN79sTRE/UGn/lzN1h5G505ddlQfqfdNLKjiNmRVGftkv
seMxDPh6L7UkHpmghRERfGwudjHSnscS6dB6B90HDq3TfIMnNmTCJLiIgkBSqboa
Ckc3hqkO/qcucoBcK4k9Uw==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=128)
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect key_block
SDTHhuXgqsjnyfqkamY8GeBYOjpZwOXw6Zh1v9Da1E6JFESgc8MzOt8ge521WiCJ
9kZtd3VAdnjUH2MUuiAjddWnq7jFvkCMlV/NeBMZ6RBDKNYN0EoQ2OrOLUc7SThb
L/lfB++CXngfQdbf5LJLsDxLD4i6FDADSDAOrDGTuWA=

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Aldec"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect key_method="rsa"
`pragma protect key_block
FaUDbdQmhmm9RqBWT7j62hCLVWsA+qf3/VHOddxuOzau5FjBlnkHgZGN4i1elEbc
OflpP7tAo2gz9Y0cDY/vZM6TgNe08pq0v9QZXLfY0CqTn6My/Y/NCsDp8F2fUlhC
+wSw6+8ImjafckeXT5jnR0HwcXdkafn/iDDf9SrmzFFwE0FD2LBWOK8WVJ4rICvp
A3LsVgHFTx2KKgs0nMp+aXRmME+hIwPKI1FbwM/rt+svBlKZMosgASl7GF8IfJGp
NJmKA6XyaGscEhAvSthIw4H5h04B0JWJDPSFNl6+mcmbNglHmdpTX2PG7qPDqpuv
LaaTgp6m3QHM3uRwCbJ3rQ==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect key_method="rsa"
`pragma protect key_block
l5naH+6J3+NGQ9q9LY6wEs0wSwgg3/pOYRWHrBR+HfjZYr4E99lybadQXhNeoi26
65CyVnsW6O9DeNA7HzWP6bln59ivezNfj+aymy40lvGtSDTlPJNcED+BzXGH97sD
Rrjy7kxs9xdVIsX608u3vXIsIXI72dtpGYiqWV10m0uKQ3nGHIHJn9UlHZK9yBwn
Q6KQZCaf+9n0JFI7hXlKhNbQehdge/qrmi27THP82IX0kKnhXSDTdA9Vo5wEvwke
wgsx9yzsjaiQEbaqZcKGA73a6qcp8XWR1o5eodrw3cRY0u/NMoFWwG0G0+m1EL7Q
/Go8oVFIMHx1rA+o3P3X+Q==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Lattice Semiconductor"
`pragma protect key_keyname="LSCC_RADIANT_1"
`pragma protect key_method="rsa"
`pragma protect key_block
Sv/lgH9+jRXNqdncDWec0Gp+IVIlycu3D8jLiXcK1bPmv87etGuNYn9sTm03fZH0
n2XWAsIyjOpWdAM3EvHe4pik9XO6N9P2yPduFyiQfhSGHsaO45Pb+476JEZMSZd9
sOZABNeG5GnqdGVfv9Y0S/3ZnKd7gj2Y2by9mBJVTEiqKBrt85RbyuZ3ee4280G3
y8ejhfJs2oKiT50uYvZTXQW/oO57ISlP6gsUSlSwezi3Lh7o4zej5AmCClxJ0ZcH
MGyWeQ43s3YvwhXGT3NeIgSXBVhBHqZ239Y+cuGawjs1hEmTpIH1y9mB127rMsso
xA9MZKCdMro7YQX2TqZIvA==

`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype="base64", line_length=64, bytes=208)
`pragma protect data_block
dGbFRfdaG2wJC44LiaLbc3INwMiPbVhO5gzo/vSXuUljkawnmimBYWuOCUd9YEM5
OOar7zjNDuQdVBi1SFhrGIQUCb3nuz9N+WeuPp00dG9tX5I/0jeQpmPjQWZYG/Gs
1iGK9FQ8EFnNauDY/gGaqQgYTVgPhUcmxHajF8lj95AmK3MsRsy7VmQvukNZD/Vy
cVa2dFmuK1A6N31YJtm4gC4yoTHIFblIGJ1gqQzLvBD7NQo5snsymLL/4E2KsPNa
lohXqHMr9Yx0dgPxZ4NaaA==

`pragma protect end_protected
endmodule



module SB_DFFNER (Q, C, E, D, R);
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Lattice Semiconductor Corporation"
`pragma protect author_info="Lattice Semiconductor Corporation"
`pragma protect encrypt_agent="Radiant encrypt_hdl"
`pragma protect encrypt_agent_info="Radiant encrypt_hdl Version 1.0"

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP15_1"
`pragma protect key_method="rsa"
`pragma protect key_block
j4uranFuSGpBhFQWFfdIPVMMk9IMddqjhcaXGzKRf7Qnt9URNVvXlkxT7epaOw3o
PWImZiVxmhuY7jgycAHDmYFghdHryUZklU2CEMvvi842BoqiT5YAQ55O++E+7BFy
e+tQiL3M0F8vsEWLDvPvO8tvYZzpivct1Fr69ICzho3iI2Snke1Loi96k4O1Q1q3
NCjMv1+c6GqDeEAuD9Ckre4sRP4f9tl9ODt5DJdYJhogDvTWYNDhXn6ZOo14b6/1
vXOAfu0Asvkv59Fukpe3q1RLdOx50Su1AeEJ+CrLCRkhHAvdPqOamHVvEVBs4i7y
O1I2Iskc2ZiTkoRIezQjmQ==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
raCmVyxIZaKm9qK9SHE+tFTpd3gOrLu+ZiIdwfR6FVTfDm77oXb/+ehkhLRt30X1
5YU1g6N4DBECQxoOg3CSzF9tP3kzRAJBoyc+TYp3JH0bKPiyInwNul+22hgcGvT8
Q47+VSpJ8wkYoxkY8wW5Sv9Aw+ZJQp/M9B82ab/6KzD9ty5nH4JOFONNTJlKw4BJ
wsKwa5Qm7IZ3Bwbb9pEKKEneMvw5RE9Igqv/nrlDjTskyM3sbByj44XnswOTFg7Z
sULTWMXcfBOgjKWeorgJLX9A6CWes7UlwD33u4XY6xKHXy7sbEAQb0Alk/GnEHBG
kZT/986MGjatrd/VbcbyBQ==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-2"
`pragma protect key_method="rsa"
`pragma protect key_block
ZtJGKN65GbSDvLr4qNm3ecd9VtWqiKnEgXA4gfWRAPyMlyk074YHnCKUGcee4bBg
Oo67xtoigt9gyu4jbpOjM/KiYEmorwlCZGI1jtyO+wR0tWcOnqhOK97fm2Bx3ZrP
HYWDKlPnyIr8WeMxhWHfRxF/PBrs849Kxp1oFi59KeVju5w67tglf0syRxQWQYcY
RAX7ADNRr39nP4iwBfRVpIXPwyt1DPqZvFZkuREtsmi2rDDAkHwSxuF43jNOk4Ok
YXp0ojKx0UoyFiKSIv1IYhee1yyOJAQG0n6q4JdskooTobB48N5lFTqEou/sPiHj
/UXrpHJej/bjyqK9xp5DQA==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=128)
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect key_block
vQFGtm+YPyYRtnOJBvjtxq8w/oqZZXuVlfg+7qJt8O6NNQd3qek8oo7m8GyLGWvD
GRZ4r4n1zjuboj+BLU3cc1+Az7WiqnZJPe0LLMXysl7kuVRQfdSaDhVianOKCqRS
qqJWkWMKuLKbRgRj9hiB9NfbfJA8CfZWy+wj3XB1p3Q=

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Aldec"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect key_method="rsa"
`pragma protect key_block
pQrqvxw8A35qT0MZZE96extG4WEQ7AE3Rf7ZUsK09oIvjsVGHnnmKxK6IScQ1Pzr
rTSWQGEQi0LqPsHOC5PubfbkAirJtdckhqaBmKIBMws3oQPmh/04m2saCBEvfUDL
Q26dIQZw3HzLWVYv40oq2r+mqGRFvGlwC+PcH5RRKU7p14flYPB3CmccS9ZaFqVt
YIIi8pXF4JdsrIkG3yrXWfW2+n5GuPB36wmByFsw02/BA17B0XG4FzRpwZQRQvke
lDKTrOmCz6L7yQ5y/1YReK9dpdZdGXvMADmgbpgcZBRa4c3kiF84U/130AkdfsOO
KZmmC6h20H77valMuzqBbg==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect key_method="rsa"
`pragma protect key_block
JByJHF0M0CkhzxJRgf+xM8Mtzkmbo0Ca98/5cuAYrXOchux5QsNpJ9+Ua1FdBMF5
DNx9p63jrQ9LkK+VDOXAswtaQRYtTJuCDToTOheWSlhwr5pHZql5jKfiqcGvBVXw
SsPFlSIrLPAvmDljKVGgiSkpKeAAXdFFiAxcFu4eEsdUOwYDY+4n/TfvMB66nF81
LkWA2y1K3KOMzLpvB98oSrVZwT95F0JhkVEMrbEnM9goCHV4R55zUtgKbJ7VT7jw
qc7fZAkbjIM9AE3lXegFDQFNxN36ZSOEas9FMCNBMNVAZ5QlUAaT5rUVdxpwzA5T
ec6qT1Miew3HFHqAgpNLyA==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Lattice Semiconductor"
`pragma protect key_keyname="LSCC_RADIANT_1"
`pragma protect key_method="rsa"
`pragma protect key_block
X8F+sktHRqtF3+D+bZ6ymbV1zHPNZPjyIj2B7ioKbst/m8M42eGiRc3skz/uZkI4
9wEQhJ7bvFuHmvxRC8nQbw9OklkbcAISGqQS1/iKqZSUbuW0ef2IOSjO7nh5CHGD
mo1HTOgWIQExepUhQviqBxtISRGP8ukDVKvBVPrdRIMrzJud9X+ECWBmEIKaLRB3
LBvjejGrEzE3w6zeJjt38M3s0a45gdPowRLFJsrpgzapqIPSnK5Dtv2BA6p5YM8J
LcGvxRyvv2PDA21Nz0EhioH3eunrq/AcAIYeCaDTctvqTApiQGx13L9tmnnM3HpS
zF0EJkunQy1532tPnx+0bg==

`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype="base64", line_length=64, bytes=208)
`pragma protect data_block
fawPcbK7a/fYA6UY9vvpF4Nf1k57umG0GQgwPfe4//Rv/fezBrCde5WBqV3jQXox
XsPSykro8nrgSj1p1ASgmnby6ybHopxsV+WlFZ+majqYsrJDV5zcMV2POLvyfGXe
ROVIT5xgLhT9knk62JTNQNksMlpysrdDkMUUtww2X1e2/XcJw6MxKj84Cj0HQz9T
xWamw32TqfaVtjsQJxD18+9GNPBYRjFpe3lxMwazRv1vgjzZenFkPY90xKvMOZIX
KFmT5ZVTb/Iu7CUxqnEvrQ==

`pragma protect end_protected
endmodule



module SB_DFFNESR (Q, C, E, D, R);
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Lattice Semiconductor Corporation"
`pragma protect author_info="Lattice Semiconductor Corporation"
`pragma protect encrypt_agent="Radiant encrypt_hdl"
`pragma protect encrypt_agent_info="Radiant encrypt_hdl Version 1.0"

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP15_1"
`pragma protect key_method="rsa"
`pragma protect key_block
oUNmrlk6nvgbnPlEAJMWtdkXVUcFYba6XvNqgKj5YDha/QK29NjBOBq1OXwVcBhZ
8uCbmz2HoxR+zCYPJucGr4Jrn1UA9tpCCKZbFYdNkw4ONqKeRbK3/F6tayMZcp0N
vvPVfu2co/cxy/E7h6AU+6PHXN6gzcchaB4DBvYM0tJsclTmmAWz80JWk+f07kyT
J4o2m0SfFANfESUBIuOYJiyeDFTWvqSQxM/c6xmB2Jh04N50/APPRhR5EiWklhmX
106QXlayHTG50HhXrdCD2qzOlt492xIl+n+egsJfJHKEP6Ygi3w0cR7I7BQmLWM0
fgiUZEFQHpYAfAVgRS21/g==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
kpxnnJHp8ndmx7G+iMHw8h76JrUzcCkHixMhL/EPaakKjDokcTVTE0eHa9VIeq9T
u+xIETfw/1yNeTub6GFC3cJeLXcz+MudjdgtclFuuGWXRBy+XVBIOCnKhfycCWdV
uZOQ17ZaefNbF7vh6BTGgQy6AHB5+8CRQujoRZ/cU/OeV+DoLFzQ1YzJ8F3lfL8N
dmw0Yb3MqxfgzN3cGhOUq6nmnumL2P4UVcxYdmcEy/+x+uxns8Ddboc+WDxBxcYi
Sxy0Uup4z4F4/PMFk8/H6ale8FKZSyAJs6ForTrgw/xItkHtgi1XY6LNp1BitiZC
RyphNHeVJXrUtwRWgH0oPA==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-2"
`pragma protect key_method="rsa"
`pragma protect key_block
Xm9nFGqFOY2V48ys50/vpj5wsK2NTQFlehvO4wRhhr4/OGQsxt2Z+0E6ztEA/S+f
FcCMk6QsD8dsDVcx3Zc5k6BAr4Hz4lzXiLJVFhRjSEpu+6DU/kNVBNoQG3rpRxas
AhQ7bXgFgkaVpC78K7YrZLIi6cA7j5t32PVw8/H+wiPBU3Wu/PojzmPN3OSBRY7z
zOlZGpkVpgm+aUZEGtDVG+ELZpvPXkh+qHhXR3W+655Ow/t76uhWup39pSRjJwho
fLg34I1zKVKHQo7J7QY2FxaygCRkaPX0DF9pwj25aL1dreSGtnNe5YhQ4zjd4zah
w7dZDBDZN6OAtP9P1cthcA==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=128)
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect key_block
fjmGOPMkubCUTJLC/4Gi3rHNL5UzeMxZlyuRAvCNqIHKVT5CggEOTXr5sr0DvXPg
Zp3hkpqA0D2Y2h1ZUQarGvEpDC2QIicdzPl1AWgRytba5Wnr2y314jk8Dtmz0QjA
wok8sQysLDIxlpOjIuEwmdZiVNLkje9fUiCiyu9GA/4=

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Aldec"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect key_method="rsa"
`pragma protect key_block
IjEy7YLNoxmE3qZDmQ7zKNhcT/0PBNmOh3MRJ+4JabQEQ7l5mthOVJ+b5Mpny65u
BSkOGJT9a3EjTdikP2hA22Mnwb63kKxihpmxZHi7pPTemtbB6yIzhXdnhA3YDi4r
WW+Oo1CiW3BOPCESG5i7yuA+28RHT9/omNK9ZWDASxAcM4d+FkqAT5HLqc386ysX
fJxbADQHJ3SCPflnQGCP4ELB5sfBXg4PHvXMUvrt7xdHJrfcdRvr/8B5xHm6A4rC
n4wBLd+QbRtoJNdIH0nyIi40R3R2G5kNpRRR98wLS4pUea4v8qsWsT//A7Dr33pz
1tCU63eHUUXewOZAccyNAQ==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect key_method="rsa"
`pragma protect key_block
GRYxOCrVW7yv8flA/fyreI37HGgO+IyQhb6pS95F7ut1t1OQ7LIp7DMHPZaNsUS9
SJc+DkpsrxZ26NWq6WNxAERvyTgFVjnTGcfU6l3CY+03sCrpKrSCnK8TqYvj/XUF
tZVBC8ablsA4XWnWAdxR6auHjDfUaAgvXPu83DzZY2ZNdgcIgMb2+/0np+rF019L
evhJX6mCVTP8RbxcP0VlVHuxMKKbky9v6hXsft56j9DrlC+bx6LTFwlNRCV1euI+
fYznbFXs5rM5goH6Q1klDMskuoW3FpCK0J3jM84reqIZXC++e4tuItSVAHW3KYjF
asyJ4Q89qr4irzVIjwJMYA==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Lattice Semiconductor"
`pragma protect key_keyname="LSCC_RADIANT_1"
`pragma protect key_method="rsa"
`pragma protect key_block
qFO4QHD7RCQv4TgGinagbEKNAJUJxy6oEGYZJ0G6UuGgcXyxdxqKd+R1hf3kYyPj
DUjeqid0UqaP6cyVT9ltc2lxR+HkR/QSoc6HxEgsaaekI6CSrgPnBlQYlHdE+7+z
Cp18t8kg14DvHc+GnSqW2SXln40EdzVdD7QX5wKae/s3d4EWR9Gi/YdeMHcvN50p
bNawZ2pzoLByCEaSLm9bPtj0Fbu17RXGIrBnWzPSiV/RZE9bdQtta/uTBxB7CxTH
zF8LuFBAL5Q2PBwsvXKPtsTisATjc3pabKCdDNOBd2ZQteslFzxCdvw5OEsPRkDX
eEvPlgVATeo0iCm455DnDg==

`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype="base64", line_length=64, bytes=224)
`pragma protect data_block
wozkx2MGGrIxcJseURmnapcTOzQWfvUDsQTxZVfXtEq3XVV2b8z1qc6zCfh3x5NR
+PKchiT3RT/6g+WO1RBT1su6O5ywuPFPUgIOvPNKb1ZZCmvQs1+BuIYU8cOVUzV8
slNeEp3c+dJH/p27RppdqUe74OTArjRdMpFNn+VGWz3hNorJVx1c/JoJnzC8LSnA
Mt0+fnxAV17A3UdNJkNKoWmv4e6fYgOq/ne2ApOkt5M+E4FvNXtGCBnbPem1LHwd
g+J+xJ/wt/jlu+HiR0ZC+JIHTKR0JSuzxiYHLdenAY8=

`pragma protect end_protected
endmodule



module SB_DFFNESS (Q, C, E, D, S);
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Lattice Semiconductor Corporation"
`pragma protect author_info="Lattice Semiconductor Corporation"
`pragma protect encrypt_agent="Radiant encrypt_hdl"
`pragma protect encrypt_agent_info="Radiant encrypt_hdl Version 1.0"

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP15_1"
`pragma protect key_method="rsa"
`pragma protect key_block
dK4FxokT48+IdNEKk2Hyin46h7syfPQYeq34cJ7ZmJqwFyiPdTAF9aLzeDXdgmdk
QHUtLB1YKEqc2Or/bN66Rgl1+sZBQmgxH8I537q9ymPWs+6UQFJf/KSrfOgYPopH
TMKkFZ/Ei37D3eO+72nul11HAdqtRGtjNnch7EJogW7h7w34KuvIOd7VC4XqFcHO
ERLKwvXZECC+zC4DSHff7vALOhTXWQwxs69kDGPEwpu49cXNInHZYJ5kIBiSnGAO
w/7xAdYwN9RIv01pY/tpbJu5PI0OD2zxOTRv3qCBdR3n1z9mLqkW8XUEvKiZm2A1
aeKofbBKldyWW6gV2fqOEA==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
DKo1RwrWrvrjKfPxLdVrfms3wyvar/0pqbWS6VQJDFJhRytkD+2X5R/CRfz1lAkk
RPVsNmeQSNO4k272UKqh0ZDLMs9aymrcg/drk/Uuex0gixay4M+7saXO6fnRsKpI
3tmhYQOb4Pz2WxuGDcfNePd1hsZxIS9zYldlg65KcZo7bFcGMCUOhoF05fWf50kU
MsA/Y6FadfgoNEv2ZNgI+g8Ai9lIEz6AbpNgzDvZy3ja0p9pBlrxfvfl2UKXe3fG
YZi3+rsmg4OxtOQZnBNr/0M8zhQJ+OFF1ZaSidqLoA6CfhKarPZt5jMGKqVtnDC+
RVpzVeeAVFqkoHGZlSwX7A==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-2"
`pragma protect key_method="rsa"
`pragma protect key_block
l8T15Zu/sbmIk2RLNxivh1UMiKW04OH1rOIWBsB+psE79nzhPvsvU3Huprwo/opH
g0hBhgvqxX0u7Iz35sUCfF5VfwwkbWeEEgf52iMYxx45Arm0Kr2Ny5DFeTA1TOKM
DL8jHC8c6dfbXCcZh0JUivGVe9ZhURtd8utHWAbtEBAscHfhNf91EwBLSIbSI8FM
56s5ghd3/NWDgOMNJlo+jzy+QhoD+jRGTuRygEvsPuae6Z3yqEcjpSTXn23zo3t7
rXEqlq3YjckBiuD4FY8vXp1Oe7tqFeFZxRXXlXPxPUuzeGCe4h2TNCIC1XGrjqlx
uaajKCNPwuxDBLaPDfLlaw==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=128)
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect key_block
EVmrxp23E9HxfKwp3gvuh1iCkKAvyq5r832QgdZ/yDmlIIOfMeU1wgH/7dFK6L1d
7yoMNYeqzOFGqjWZzIMiMaRuSeqUCAidjrr7RQ9hb5vLlK4iEqd5VXmVVPvpTYx4
CSf2tBeWxReUVmu2nyA0FEuouD6GUnqYkYxQSbzkThg=

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Aldec"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect key_method="rsa"
`pragma protect key_block
yotljJnKLLoXFeTJQuhu8wh/gV2vJkhS5O2K89Aw+ENxwIk/6K3PMpDEZ1nVcnMx
Ik4ruUK5SYwmVzMIL9dRFsCRo1LheBnNDdni0rJJJVsqs0AKqLYGLuC7R9srOz98
g2lCf1gGGF5LJ0WJo6tz67Jv65yqPdixtzgv1xX9Wct6dopXLYGQkqlboiRd/0W2
I+56KamumNbP3afXz9lLBWPZ74Cqmo82v0HeOgX/3qx/XruLV+vZRPoRBFFxEgRv
cyFEcezEzttRD3xZG/sAtFVd0ECg/Du1G2k/uruvOyRgWVpoblI4dN6bSENRCSVU
vID5KuIRKT+Z8oqU9gkLJA==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect key_method="rsa"
`pragma protect key_block
hIcnqDUQdJdaMBOAfcLjiTGUj/+HFpaCyPR1qFybBcCwCHZhT1g78jlHdjheV0J8
xM8yDRRJyGo/k+PWfbhYlW36Dox2nkIixCaWn+AXGhSWBKBUHveM1D0vRfKVoKcj
kJSBtq04jzNikpoUzYctwvuTxrGcpaInEa+JDukorz/iWxotzDZqwA2NW7WjofTt
yV7RRKMh3hbPsJ7RrLWfV5bRfjNxoyxFV30/zr6lUMdUkf0yH7nukyeiHTqN8PYM
qyeivrMaxgF0WHhGCOSdfMV2Myz1GzZ0UYZFR/X3GPJd6+gApXFecehvExQf0DHY
baoFMD+cieOGH2zoxX2Wbw==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Lattice Semiconductor"
`pragma protect key_keyname="LSCC_RADIANT_1"
`pragma protect key_method="rsa"
`pragma protect key_block
QbETc6WZCXEZQ3otWZvWJRMR4CagSjymsu7jADvCy27AeAVosUnJVnUMiLpYtx4b
BxtQDMAYx/F9I73fXQTl+FiSqjsG4Sf4ScXR81qV4cH9WzPHub5/eg5x3Sy1uY/J
IXYMJ/aNkNdZZ/mCO18G0QcUjmz+7DVlFJxkXbgrA+ga1toQQH6ALBnjBujQFFQo
/2QgRm91FfKhAfhTOv26MWfy+X2Smj0MDcjavuUui8feeMlpKT3LJHE52r4bBipA
sH574g7RTesyeGORKc1SmnEv/3SWgVWgyhsyPsyagTQhvEeoIoOR1ED7y6uqHiVY
OFKP9W2g37in+t9xYDVSLQ==

`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype="base64", line_length=64, bytes=208)
`pragma protect data_block
DBn1DhfB0i64RSPXbSsbtiK0KTlx2rTSr+K2EqtLwDh6qmSlABGKOqCNA9kn/pqr
ZqQrrQGvmkVGvwNNzbxTNbLvZwydWJzhaC6i+JsHA+8SzfykNE6q8E+QxTThbATa
s+IbLE5amFZtn6y+kol21+DY3fageCQPT4e3jt9M51NboWla3pdB0MByUS9+qtnc
eOP4DJVzXjy/Wwv2Q3IGJz2B8lpCyvLeip8WBbcWVkdra8eFnxPlWBbvrn/txPqi
qfEhDCTZ2lIC4syn+cDoRA==

`pragma protect end_protected
endmodule



module SB_DFFNES (Q, C, E, D, S);
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Lattice Semiconductor Corporation"
`pragma protect author_info="Lattice Semiconductor Corporation"
`pragma protect encrypt_agent="Radiant encrypt_hdl"
`pragma protect encrypt_agent_info="Radiant encrypt_hdl Version 1.0"

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP15_1"
`pragma protect key_method="rsa"
`pragma protect key_block
y3WX/WLrfOESIzQeNnAP+Vmq2V50Glqn05tGXn9NU4bOmzxVZURFkczu+3DmcveR
RYEfglQersjajZQWVeVnU1NiXMgzDVEWkLzWYcwCiVpq/tFFkOBuadY22eS26Tca
6HDu3gTHUed2yBn/TAw1oT+wZpzpsPolujV/zEavOFNEMB+Hcpf40YzjoOOtXhy8
P/ClZYoXd0zkH7cImPp1VX4OI60mN9RXTvyXk7e3BZ9PTnrp8uUWUXTxYVB8/7h3
s0G58lpAri3JlipMWkTzHlz5wLDKJCQPpQnryZ6ersVIPp1BMa9C3WGPuRWvWFIg
fpQy3/qiC3D9JuS1h3MYEQ==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
ge6q6MuH5AaFOrKLzcPX1kPgW6K3oWAgzIbJbrWtwJ8Dg1RsmVUFiYzUP6gNJuGp
bBAWMZLBvSxz6U5dDUvasrd7ouQwJxmVmnXthAwLbK0Xeeo5ztQUAJG2C0vb/ATK
YwcUIPnEWFwArmFF3+eTvEk0lPpFd2D8Dk5EUv1i6fkcRNBaeTMwO4JoLCDfpSJs
wobopJsUcfM0m91vSq10XczSloYnfnlQv1v/IP0qifcRGfiUEQaB16+3upNciRWe
e77v6IYB2q9A8kOeOqfg/No7d9MgW6V32AcJ+55hg0PQQJPg4CTOuwPDZRhrVC6B
s3fJpvh+MqMkqJuHxkgApA==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-2"
`pragma protect key_method="rsa"
`pragma protect key_block
OiizXzuye8nD86MJXQXC7YUxkv5gQQqbfHMC6/hdRcp7GKmYa27z4dIPUZn7pvg6
NpC7l+KKySFHYcYiAA43y20x/C8HE47vP/mxxtllW3i2P/peMtgenwOS3Ywj9hie
RK/ztfvTCxy5kXpAB+XpTxwZlLvRQdzNtHN4Ko7lYC1DxcBGA28nMXbE6rYl6zCb
IIpNj1C3W6IYLi9wcD4I0ivSipJf0ttoN95NUsttSaIBNcufQIzjKzJDQWKfZw6n
VBG+sx84VaETpa1YhRXw9035WyF5U2RpRibHqR58nPM9rWhwkhJKHdVfCqzECVuM
vvXXqHxwT8XfmOFPjsGW4g==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=128)
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect key_block
jHd7dtxpMgZrfuOorOPNPg3b/gnwdE3sPdDwC5nwumajLZlRLnb/lyS9D0CXo6aJ
FPsPWWCuAVNiBtr1koTOG4kkLPR8n7hNMS1lRP54oqvNEmXTxnl7+f0qJH2ibIVd
EXyabOIJNis+GLHeoONgsdARwyM+xYe7pwkrD6TiIww=

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Aldec"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect key_method="rsa"
`pragma protect key_block
NfR4wn8ajcUo5zvCQdmkWzA778oe0Xj2BaqfyVqxbBGjFL6hSP714aLwnvwbKMzp
TgWqh7juVLSWB2gkiaTr4Q6NnJ9GG2lm0uCqsyWyY4lDs26mJ8IdOy1VF7ud2wms
CHjIybmoZLJ0h4N3EKQGdo8E1Z4Y0rjcQMaiO7CyKgar/cQlDbl/sYm/x/FkUF5L
YMFBffFYCz8tRz3zyn+Qgl6TqOH68/ivugn4dLZSB+tmqWu8BWiIzoq3IAzpVTJy
o1SI5dd2IfByMxZw5Oyr1h3B8DyphQGEYrwxBs/6I2BFlE0dBHBmFCkH+nDV3hmu
pZWoJNonTnWcLSEcDuCT0g==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect key_method="rsa"
`pragma protect key_block
aUJjTsY1PEu/RtagFMpRYnAqa5tB3Yc6B3mftAWzd+UYm4kLgQg6vvRn4RDc1hFp
XKYeAVN6l40E9EVLdZ5hl0evJ5BMuhOHHOl2WhSr1qg/kiogrYPRgEe4yhAd4FFY
xf0H36srjLcNbY3XWLAFtzU83D48sa19f+hKgmECqd+xB3+9dg65LPYtghqZPWA2
+APBu4q/yZ185Ft8y/4C+ZpUsdJod90125j9VL0MRdX+ApaOFpPmTpaV36Sg4K0z
AWev4hmkfGzdb2DCwzpAxRLOOpaedqT/7PHnyuHLJGu1d+EVGI3uayvc7merz9xv
E4kD3evzu7ziq+ldLUs8YA==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Lattice Semiconductor"
`pragma protect key_keyname="LSCC_RADIANT_1"
`pragma protect key_method="rsa"
`pragma protect key_block
uo14U0zbrgXU9mduCbt6BNTMfi7lp8z9Y0n863dTTFKq+uGbXVw9AUyVhAIGIDgA
tHl96xZ8Zj51ZYnM6GpAhLtI70hRGLtbSfn8vds2ygDjW4aWskfmuj88IUQyxI6w
JGrNVMe2KpgkthMawVz0V7V2To9TuqNYFAmoqNTKYmsQHQqlWfRIPjMc46iaoxpa
c7Xv7SsvPaXas0V+P8ZgLerGOgJAplBqg3pjPTts/edHUQXe7vTkJPHOU6lVUJIX
bKCPT3DkYJtEsVniJz5mU46JR+RqfFcAYrapwGagdqYtKeLxdYtdu7vYvD00hF2O
HKobQFHjx3Xycdur+yBFEw==

`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype="base64", line_length=64, bytes=208)
`pragma protect data_block
dAtqqxwf/XqGu3FV71zBiCioXimEzXq+vy5G4htwWP5c+6pvN4ILYTAKbyXFcXC8
G6XxnVAnAyw/QV65VtZczKww22pk3k1+lh7g8fRdt30xuxw2WJHjJeFn8kvgSzc2
dVA8cx4qzza4UonNszLePZeNHtcWGF+I2Xudx7xyoEjwgoRBwO6MdqsL56czlNsm
mCZajdR09MIH7lz/4UsZ4p2lvECpqQgPsZnbMcrFLG4Mpp8ujA1pX2GKu6xp/gae
HhDmO5fdq7jog9oebh7VHw==

`pragma protect end_protected
endmodule



module SB_DFFNE (Q, C, E, D);
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Lattice Semiconductor Corporation"
`pragma protect author_info="Lattice Semiconductor Corporation"
`pragma protect encrypt_agent="Radiant encrypt_hdl"
`pragma protect encrypt_agent_info="Radiant encrypt_hdl Version 1.0"

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP15_1"
`pragma protect key_method="rsa"
`pragma protect key_block
XoCP7981tHvJhi1OF5wkNGEFJ+KUza8CMScKSoQmkocYSsKZPXjBuyXkYsFa+ThY
RA6XtpnmnnqieI7LdxlIo4ndze1W3VblSxEHxoLxbjKNkqArwVcwkzTP8RoZveSo
8KAZZb0lhDAhOgmfrVF+ZM3CP1ejdoFbMFzCa2cIOQHW5GdlZY5GplvM5GNDJQOG
s1cN4zcFyc0jL06/+NPqbeFTrxFsa44iH+PaWHdIcDzXf/HQDxp2y5GvHbr3CqtE
lm6tfv7Mrm0x5qC/XTLbI8o5DUfEIfXvACLDCb6dnRvIxLJforNOOEUn9bv3SY0K
rDePtq/jc9OV7CE/cvU2tg==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
nlWXQJf0FnfA713laDEd6BiLkWn5T3pbqxRkwm02XdL5QlURpLV5aWJ32hhZQrep
ezkLnBQvag1GCSeFljgFWhkaygDlQuMYrfSUin4ehydOEnEFYcM0pMxMOwR5P/0A
cosnI7SXhpZxoQOwlgR/RCHAiGxPv4o7kI+jBTn+6SHaTojojZ6ZMa7AcYCuOVvS
uyeBOOiHYN527Hx2ElBHbjsUmX5AHTDzDjUQdiyD9AzW+U5XNJIUF+Fj96j/2h1X
jXRoX1zQDf/4qDWIw2SUWKIy+UZBOAtJIPrb0rCBOnh5eucH4jImwpfNp7X9n7NF
B1s3/BPWJQwVMC5Yvu99Kw==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-2"
`pragma protect key_method="rsa"
`pragma protect key_block
ozz+IscLEMn9UxTBotbXnkbA6vuvOv1YtbMmGhEqpAo2JYJMf0Dbvg3cEVY7APFd
+/cMy+INjNy7UAKw1tIqo5SVq6CcoAD0NinTAwdUcSHOGp21MS+m9XUdq0yMuuIS
T8tvcuRxF//fLJMfSYZAdYThKE6dLNsfuJfbfkSQzCpIL1YZM2II7hXcJjLoIa9j
orAfBr82f732CwUENvcwtAhGdoyMPM05MjCet0yaFmHLnGwemAmvFLj/KddIKzbV
rSmW/jbyu842oqAfLKYXBgra6BhrOCtQCaez8wqZcW3xA3FI4JaQXDbdm+mluvDK
O5rNWjhm42F4J5pvLlM+gw==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=128)
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect key_block
qwH5DnF3lntFP/d/iKQyboDZ43z4YFjSGiwMPSAMzcq9OynPYH7Pf4ctaMU7ycjw
BKuBUxBE9mpMmOv4+qMbrq7era4L+ca32ZhAGMGDwlPGVK9v5NRqxZ4K+yQ8xbYh
SwVtj4CgrZJ0DCNSjZIr2rS4bBC5kXzv369rnHmQa4M=

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Aldec"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect key_method="rsa"
`pragma protect key_block
vYCj6YwhA00LooyMF0bqCA2DqiKC81HCHlkgXoQtUlk0IO/7kEUIo+bcNGAYWdbY
xBTTe+32YM8o0ftniM8qUwAGF0O9DEsCig/r0ACLHIskw11JPJNHL/UVag4IyMdx
UemUrTtTv00qR1oLviI+tQlOCraTgGg/9TzN2dHApDTaLMKx+ZoBEiM9LDjh5ieP
RUy6a6M/fY5ppoWBTu+OQdLZtm4ZOb0npEUktqFuwjcvBheVH6MY/cyPrpKy71my
bRdCRb4L3mMHIqBVwsUfVPbiz8UyxAMyXECaFh9twaFAUrRzQsFMD1RRqLXk1QES
nwm0bQ3lcDr+3BXTimiiDg==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect key_method="rsa"
`pragma protect key_block
oHEDy75HqDjYMrG2PAoVIQ3o3j44kFVJRS9bTm1d2/ReAxtkvpU8MoERKrRd5BoA
nPBfRUKo98UZ/HvLtwVKcwcHAVMhdy8Kex/s0SjgyvGXjRoJfuRqGJ8fj8Y5ZqRF
+FAlbOn852aZT4KQ5yZbRYamo4MgMDPIGLLqvuWn0vFT6tfrFK5WBUjhBeV9vdr8
EEp4ajlHzn3dFHroUfIBm7NPZYeUy/FHcc5oLQJdLSlvJxTFqm3TvoELFrmZU5g+
jwTsTRAM7skwTd7q9bPRqEBQUXMSbF0taTccwus6pW98tNPf2EKscGBktlHj7oQA
bs+pZL+t5KzcZRBTJGQW2Q==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Lattice Semiconductor"
`pragma protect key_keyname="LSCC_RADIANT_1"
`pragma protect key_method="rsa"
`pragma protect key_block
qFH4IvUixFBWNrANOdA/a0Q8ftk6sjBpS8M4vasbiiIjz0deghz2EBOI6zjURmis
O/os9d7OWLJs+dWhKhDU+N2n5qGZGdLLTK3CPh0yOsDU9MWycV/619vT1qEgVtMt
51x5aU5k7QB7XUrqCA0MEFkAtAIEx0cF9t98b7hYyR1VcJ+Rm3PpVNLJLweHhwmo
HENBTw1IwGqKIsvxwoBHpxa8k3D9eowgBbHKWbFhcTXgYcj1q4VjYxjrQC62kAIz
N/HpKsy5Efj2syYgxwWIJA8XqZm8vLW1kMZG5ADBz9MWVBwzs1b2fecU3Hd8CWaw
tqg9k6IZgpKifzYGQlRWGA==

`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype="base64", line_length=64, bytes=240)
`pragma protect data_block
TcCY8cjljU5QijIuuhS8Nsra7eQ59eAZYsQMNy9uCeM0GMMAhRrrPha8T4iOQTRV
1aYvAmlTMFOwsCYcL2i0qVBppIDotj2tVyCSBskvIXw3wcsCUMQVtwGbIO9r5U2q
beI36KVm/o2B2j5395oGC03mmHZY0ZZPbQVYOnCkfl26652MAdPASQnwyEyDHTH+
U6mSBBZSUnlRf+cM3nIm22jWTnS60/5PtenohApoYzkny+YHk731MCJ4z+a4o97Z
cbApdqtGQtcuDWa5zR8qUthfSGUTGVRYNEnTYmUxyAZnqiTemLV26DHD4jPoII+j

`pragma protect end_protected
endmodule



module SB_DFFNR (Q, C, D, R);
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Lattice Semiconductor Corporation"
`pragma protect author_info="Lattice Semiconductor Corporation"
`pragma protect encrypt_agent="Radiant encrypt_hdl"
`pragma protect encrypt_agent_info="Radiant encrypt_hdl Version 1.0"

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP15_1"
`pragma protect key_method="rsa"
`pragma protect key_block
mPbu6NFCXiL4j6S7vFhzqPFsEVUkt0TjQHh+XDSJ0RtLI4PFuNMKFe+rohnk3KfP
xOMhkWLXdG9aB1xT5tFggQBxgmj5sybOSlkbLGJihuzCMumaPNbsIHrsekAwy/gT
nZq6wFnPYg7tk80puz2PVAz5R9zjnE06aW6Rbqfnt97X5Md0FSxTuGAK3nT9oNuu
FeCsd1yM78o4Mwkc6MSy3nxV1HNFNq/kcdETkZ5aR7NT4rqFmNVVZ+VcTc2NNoY1
h7NoxE9jGl95Tw8In6KGWwu4+71rsmaNDoXhKNEbqTWPfu+4JYR/AlAqKdwbAI8Y
Mo7sBrdA/jWFlHyk2cdXHA==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
U7+LnYoIRqmCWA64IEOOG8yPXn0a+hNPSy3GD3NMnq+z/MB8tGvG0WapHCz0EmXP
okx3dQF/7g5OTrCs8i0aEsdb1qJjDGuVfP91+t820CFQVpAqpNwm/kdoMz7kHAZt
J7qR46fruaYKeBCKACg2FbSoNEL17ed4PTbz7QbHqHH7KB8N7mXKTRrKxttzxFcE
rU9SDWvDKZ22T+Fi/7p1Y8DTcvVlaGFBDC8CMWwMJHaOVrrH+GSgYj64dFCKL/pJ
DNX7EoaJ6swXyAf5j0mbbk3t66M3inYoPR/TM/XsCJotgfPQsKRe0Exm5eC5Dw3W
ez4aVrFWtTUQ5VjebPV0EA==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-2"
`pragma protect key_method="rsa"
`pragma protect key_block
af6pGueNg1Z+quaSrDvgQZcTHv1ssRRKQZzqx+gfVExrnbRjqPUWmTJZsSSOfLXV
XeqA4rt/OIxgw2+qD+g6DVZvJY17ImFZ65W1xAMJIG71q66W1cIpR7ZZt1qFzoEq
8BDfy1+sCK4fRwnh4SlAW3pojGaCHbFZ88/v4oOvRWai8eSnk8++TE2gFXkY8juS
nD1hnspo/AOcjMSppCzV6yEdLfFlqMaZUuSfI7jddAdSqnxjbJijj/shz2i1wozJ
2Zy6apaKdo/IvYIu6nO4+gru0PZY2F5iiuqWutveZMnBflYS/biAn1aVuyMdR34R
94Pee28Neji6xeGUUuZvNA==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=128)
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect key_block
Jx9CBi/tbKjj3zjbQ+MDmWKuv0Jy+wJMrhUi5bZu+fCme1RI3CCjfOlFL+XK5mPN
rVq4X+ldzKwKluBL0MZk7ukSgt1V//8bv6aTYwVyAybHDDnO5uUqOfUfpKvrNHMW
HZSvqnWlcxpCI/XwK2aFJv9pHBayhw5nbJ3gUUaNFvM=

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Aldec"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect key_method="rsa"
`pragma protect key_block
zX1/kYv0e/2h0bawEohiB3u1hSdZvJazldi67r0kGNMSJfXS863gXflYBAtNxH+/
hdy18l7jpi59o1bcQGlC6RjX1NIbXRNakePr+lp7Xv7r2TRmScEFMTGfIqCu43Bl
Mk3DW6ne9/xXVlr/sBYVr+y2UN6t93lDgZT6X4hOmgbpUAOPWUsyjo1k7covVUVr
mLMP7l5wYlsLeJx46lVOqqiQ2UMaxoj/GUAyg4Hdtdu2AlrvTELz1M8GutukbYzb
spHcHR6AaxLHyWeQW/sqWcyyp/GrTIqKKLZgMIxkccKshr1SAUdz41iKMfRyH9Dq
h76dKTeZXolLKdAVuXMiyg==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect key_method="rsa"
`pragma protect key_block
Y319oKdMudh4ctViZBifLE7iAiOdOEiRADM12xB0TV3LEv7iEFGc4hKyslVJb+Vl
FJx5dSwvIL7oeD9aU+d3lA0ZCKIsC4KwxJky33b9LtiMco/2agN8SFw9pPV1ox+l
t8ill8P6JvSOi5qWPHIOMQ52fUCEj8X4z6LtwiUMHaSga5XnQY777gwe4/1yEiaP
KNI5x1rbNLkUFJz4Xz8zOz+mhxkdUKhw8c0/tpJ04DJWtrcPTbOJx4ZW21PnTpK0
7dRX4457GmXWoYsmhbTiSrZpQJ+NpZIwxEKbenhFkO6msXbsldK37QeQ3WzSd2qz
jLiEfQl3hEfWqfUrkEZ8Bw==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Lattice Semiconductor"
`pragma protect key_keyname="LSCC_RADIANT_1"
`pragma protect key_method="rsa"
`pragma protect key_block
Qye9IZosJigCD0R5mTgbebPDDZC8Uma+LutNA1IdKEquMQnvnsJ8V8jTZiIs4pAy
QcGK4+xJV6vUGEd3VOlOHEKWrdY2ZlI4SuYJieZZ/OjDKQI+OUAzeMZYveDSMygz
ADWwmKAmeCz/rcrwNe/XFIyKkVMibqYi4XmjjCgJyFwgeUsthkUFL93N/bWVtTDR
6f04DREOSqA5nyECCr6S9jQ+Quw4v4YCC2Lp9NXJjLjfD7a0aFN8P/zqUlQqJzt8
wTWPe0W6G/dm5Tr2LwDYSgzR1wO/gVva2uGmkA9AYowqGXjidN1Tdu6KMw3Mr9aL
D9tGl2B4YHGO6u9BLX/IFA==

`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype="base64", line_length=64, bytes=240)
`pragma protect data_block
WxP2MB+7KBUH2G6t+ridyjwf3sxNWaP/89TcvtJJb1usxikoB+Lfn5Pouee2LICx
vlXzOBSHWPwSK8y5KaZQkiSV3s6lxwZxqd780Jgy0b/dOpAXxjYsyysekElH7ZrC
I+Z3qI3VFY+h9vd0Vlg3pnUd+ry2hQU75TfkZeQzyahPRypwkDlzhTEUfhbljGhf
JN24VCk8muuzwDlE3gwoAdBb9xb0D9h605RfqYjM2RF3Bcd95HKo97cFU/WeAPzw
UhGM3YjOtPRrHrDPFHfi9GYkSz/URv9svIHp3WCnRZpA0gjQHoSPZCoAce6E9chz

`pragma protect end_protected
endmodule



module SB_DFFNSR (Q, C, D, R);
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Lattice Semiconductor Corporation"
`pragma protect author_info="Lattice Semiconductor Corporation"
`pragma protect encrypt_agent="Radiant encrypt_hdl"
`pragma protect encrypt_agent_info="Radiant encrypt_hdl Version 1.0"

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP15_1"
`pragma protect key_method="rsa"
`pragma protect key_block
aBqMAh5aHuR5UWXZTnVBbqKwuFLtC8hY4cLSzrIMYiJbfNVnJpDcctORjiXqywVg
dIRalVLJyKzQkklSOKHvNbVyPyq8x4yo6TL6GURnfwI8rxhGqtokn+UPCB5fB5IU
FGNCp6T+LJ+Ge1J14hK8eYcdbg7O8OFn0/wi/tIqROHYGQzELYmYsl1c6VPLxCsk
Au7Z+NjYEeF6IRjpWNS1FkzJifi04psMB8ro++YyqMy96OHiL3aVqQazZVNQex1C
RIk1uqYRXG6i8iHxPSehQdsuckFf5VmKYL+OB3rf8yVqg3WeQO0Q/Y2yYzhcsmb2
ZNHqPJTX3adN6ay38cIuGg==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
Ybasgn2PbcAdHtTn6TmaBqOu/ZZPhqg4vylIvNET0EIEHl4+oYcYSjYhDYvnBav7
EuY3kFN2fKMwM6HYdU5xvLbjrivOap5QBbn9sMT7aHGEEdXnL97xGXqtQG7jwkGq
exo6gP/Z66Pd6ZDAJ6iw8B/Yx79zLkkn6/2evJN3FIHqwhaUJYlW5wN/hpLfIjvv
1snaBcxNjKATiTY6sTMGPMRD/vQk6p8ys/6le3r8Qhnf+AQXHLOCGwaT8AJd4wAi
Q32pQDTIhWXiXpGY7vAYWlUoCsqF/iK99eaPPPFHLJtlMrU2Sy7fXZUejduM3+Y8
VMwYEbwbXRbQ20iSCl2Fjw==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-2"
`pragma protect key_method="rsa"
`pragma protect key_block
Szn5SrmH+laOKiNAIZLGdJamhLgQywxF6c3hHiZBpF8mAyuE+tWrec/jk8QVohWs
FqDp8yAMdQyHTKSgMP25jCINCuJMKSXk/Q7NF7h1pvQMoxtn2Q+BOhyla7DmADNY
fN6dSiV/esoBdT54NSBSmuq1oaIkc7yAAGZ4YQnI94GSY30P9phVmsuIE8GgUefk
I9fiInU5qpTxc9CL13hU2i3r2TQW+uYBNdP4eSkwH40MC0BlAokz+2L+BfB1ylqs
WUPhv1+lABsurOSoVaHfk0bZJKsBIYL4EdEHma4rIBAVQIis/7dpyjW6eKkC81EV
DOfIugquvS0KAFT8OnqxSg==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=128)
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect key_block
02YJ0Zt5davORQjJr3TSGCPY7zBnU0CYHFFbnTZZwbuo2axzfmocfwYGNdSLMgxQ
2H9YHowDj3iEULmap8g4WFXwfbXIzNOav/33wv2od0SP5w1OF3x1oSNwTFuKsrbQ
sxx0NPxwJ7FEk++RA3Vk2paVi+nKMz9sLdBaAg+MEnA=

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Aldec"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect key_method="rsa"
`pragma protect key_block
agcfFUx+kqIQtv4SF/x/t5R3JaDfyX5pFx8O4fmER1VOXGACvVcSsW72xu2SHegk
p7tvFFkn3b1DxABFiZ6MxGZSCufwZiIBMlDw+lbuWPgaw+l7XPu1EbKGJw05NrIc
10H/GWMrGsn2oy2uSJwcbsADrTQgecTAzz9cdILre0nZDkUUF0Yuw3/c4NLkBv7a
v9/XuQ20chIiqBVbyM5NNuBcWVscI3WCbIVOALfHsK78f3KwHQCQhKcxNi4qR33Z
JsAvMzUvjRga1H4AOknt3iI6rpon9BK3SLxB8hZ0W268jjZqn7LWw5jHpnTN7g1Q
4kQzEzsQU0o9/jUp9FvU6w==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect key_method="rsa"
`pragma protect key_block
dN/JOM7Oi2X9X1ty9Da5/IAFeq0dh+wTfsCoynCSPtpdQ8jG260C/hr1BMsodJud
EPzm9gpFKzvR4hZRlfcugR9goGILjdPpjSJRrdYPinnzSF1RKI5BBDDwRKymkcgu
dyZw78TB65/W58o1m/hGwcazfxda9hE6ceqQyBzh6buoq/sCnzSzv6uTHLI2z83h
cy6shSHWkEJd0laMv6bOHa/GAGGwLlDBx1EOIpl9yabZV3HYkwSEWW+u4HAbz7zN
mNH/Nfpn//lxyBVRbKXW9jCNRuNuM+xWGJyyZBKAjd1iytnSS2r22IbTKulvY3ah
jrKY8oniuPe19q5QsqKpFw==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Lattice Semiconductor"
`pragma protect key_keyname="LSCC_RADIANT_1"
`pragma protect key_method="rsa"
`pragma protect key_block
DlB4yfm4XX9TdpszHGxcQP0E9QvHFGHXQ63uosa7UoZKFcp+ALKzAM+alN6uoL9k
Z4FBcLGLF8lW20Rb0z9E7cMBtn9h54jh0oqq0vCdm0SFdCh5lAGfHs1rUDEoIl/W
lM9ROwOQuThGSlZj8XlylNRJ8fDqRUkh+bf9bvXjqv5LFWaaN7fXG8uHuKohKlY0
CvZVwZ3gHkrbA5jMh60zHqjdto4dxmSNfpdKfe/ix0NgJRhS1EliHGmrQxidybTR
a6L+RxDAWJbemTXuJHaPg57URcK9mRmchbqOHnBQAXZm1p6TZObuTcTgKyCMPnHJ
e5gBqb9Ml5ANKJO+y943EQ==

`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype="base64", line_length=64, bytes=240)
`pragma protect data_block
3XsZEMsze/J02ku1CQwbBtz9m74+YfYbRLZwWyXgHdBScNI/14+eY7Ic+TEIN8FQ
LeXwIEzIbwfWn3f4x7s0XXMyN7kIIf43nfE0MpFKOag2oWitP7kw6jEBxgZ5xevk
eKxhdTdoXpJor1nTMMTXjYtukrUuVPVQmadq3o4Xilzifvd6qtSHqMlMkoI92OIx
dlBla7RMmzcdOvYNLC2XwJ/FKEtFHZHSJmT3GI0IEvxFvI2miVwFLaofPPw+XTcR
NQRLuVWeH5n3sK+62uZHdbEk1fOXoIRt8op1X2vJi6+++oGQSZ/NGEwiZW1GTbib

`pragma protect end_protected
endmodule



module SB_DFFNSS (Q, C, D, S);
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Lattice Semiconductor Corporation"
`pragma protect author_info="Lattice Semiconductor Corporation"
`pragma protect encrypt_agent="Radiant encrypt_hdl"
`pragma protect encrypt_agent_info="Radiant encrypt_hdl Version 1.0"

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP15_1"
`pragma protect key_method="rsa"
`pragma protect key_block
Q8iI/NV9zu/xphLwKy44RhxJ1bG3QRYhQROHYLuDhaIHBHnoA4931q4mNFU+QNTL
bYXHpNFy+VeqKTYBIhchAoRp4XVaEwn+36MTLAxGOZphSH6tyoyIkxeqVcLjBqXc
QBrplkuVzr+HxGuALEuoo15fT94Pd8QMukxPHp2xKr1aCY2J2+vKqrU1YgeP1MCF
JRqQz22mVuzh54+E8azbRTgT6zvgM5o3OtLKhU3IxxsMPMusULwbQqWOMsTq/ou0
RaPSm2FzZFkBZixa7mvoE+tl5zAOHP43FQshsYSVK4ALYQNFymEQVhClxPfdA4Ji
gI7hpeS8Bj3DPwfpErxXxw==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
bKFwZK7rhk8cEBcljxJWB0D2nCPV0Udx5VMMm8dilmbXVn0qh5nKkJDoEW2Eafbd
LIVnMwl2juzUxI0kSKgGrXKfsq5YI1wRjJfA+tkdtSNXsvGMQEk7V9tNrr45XpCJ
7v+DnX5H6nFXH5xZkoiCUNL46Co0NwEQJwYqB1AC3ADwTMQtobBLPTWEXQjLLSXI
L/Zmkjra3ZZFdtR2P8zaG10wd76yN9GihQ+4S0oS0j/Nu998VG145YevVMpIVvkl
bFWacpwfmIkc1FwdTtYHtpkuEUWE4xU9utwFTdGd31AqCed+CrEDk11OBgXoQ3Nr
tfk44SA5Eh+DV8JKD2Qt3Q==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-2"
`pragma protect key_method="rsa"
`pragma protect key_block
nmJHLT+QTmTUFnTaFBb7vHs11Z5C4wBewXaQEELB0xxpksqVskEDPKNS36umeCGe
0t52Po1OMeSo45R7AbbNvsPxbskYo5tE/V4jybjC77BvDEAJ++6iaBz2tH85BZHQ
FhLKxMkXgKu0GMaSCgKWvv2ybrrOIGvikIC2vQUIM5GWr95qJxkeDjcEy5t26Uul
RIoxyHvvDZfTinr+InoLuWKJaU8xnbVRcKDFCVP9ruJretACqTx+9PwrBRWy8IuZ
NNFTNCs82KgmFskoJZhb33qVWPn5DdsscqTst3WG+3d2psD1u9HInWcnBqny+PHa
3pZO75xsAQ0nLdvhytY9Zg==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=128)
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect key_block
eTngrBSAtjYhqg0AxYn9Ae3Ca8bfY3kgeOgDIl2pyif6y0g+Fck5c2msKghmty5o
e96v2qi0Sh3ApKiJSl+YaoTrqzxdfIPMYOXrKLCc6VuXn3JiJThuwcrK+csjNcOO
n7ZaMGfK98WxBYASuXKHZ2h0D67v4cYei1KNlpLzlKI=

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Aldec"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect key_method="rsa"
`pragma protect key_block
ioN8EjfiPgufPjfP3/CA/Q9KBeX0QsUCQjXcbuWci2wNlXyEOkYIAVOnCXlr/+ym
Ev0qxWyytDnMHUVpGYqn+CEZhlHYDgSzBqDG0H8AuS71u4ft1bHrjft8Uz3kizjC
ErDa+Gjw5gaYuJYR4GKL7cy21RsjYcqdBg9KXq8TJRLjej9R4/tEB62oePCGwOkh
AOifgLNJWLiutYPPByFE2M4EHLQTD/exBYp9e2E5gb53UZwVvYGQ4S4tgEWOF/F4
wVRiHtBaF1b1JSiDwQwON2AdJBtBdLDpt5Wqi9/d0cIPQWI2MnX7LxI+mtMMs2LE
oSGadXoTQ/xJyRd9vQrcrQ==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect key_method="rsa"
`pragma protect key_block
KMsDq03PFVxH4lfBt9EsxxvibIWgfFTDdk4qiJfoHA815trADGqx/WYnpIXKozCo
QmHkyAs1Yq8A//2wct9m3wjk6ZB27vj8CZX/kum2dLar9A0OK6CNnMXOiHRVzGQJ
/7QE/DbxukLVaxxavoBoxV/GXrDXELblxV0ZBhPpr8JzdYF7bKssimqi/keSORQ/
XMiBGJSda8lzD0ah1/4r01MPuJOIYCZxfRA16ZcJg9p8fdXnu4fiRaclpvoK2bVu
Y8Tet5I7EGG6JdjrI6nUwfkns5aHuGXsswtmoJzp2lShZGfSNX7KpdhoKJ05DIEe
d6Q0DD4RtG8FCLxvQy43zg==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Lattice Semiconductor"
`pragma protect key_keyname="LSCC_RADIANT_1"
`pragma protect key_method="rsa"
`pragma protect key_block
r8J2yrTdo4Jw/p32dRXwis5r50AeTR84gMmuy285CK6IBclPxExxhXYivURjjVfn
aN9+HhhQAFBCkS4PYjpr4Re64pqK3yXxUOLKFwb6YoNRmFQ2psxmrYDLEsPsZFyd
JUxtSN7Liz9SzgPKPm1r5j8AFxbQ8+GPqvXf4Hql+z1oxj1wJLCAcaHZqSe/DXrb
vZpqsnDC41Wdl5BOhPdXuqcnXNwi+y1KhDHzkNkTgF9i2+AZgypojiBUejv7ggNU
ZNokHpL7DqnwtnqdpHOV4vFoklq0Y4xncEx+mZ+/V9IFsVczRSTzY/i4okaMa2iX
ViiZLhOAYy11TyWXPDX1lg==

`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype="base64", line_length=64, bytes=240)
`pragma protect data_block
mmbexPqvkcZCZHdfKvpnt3XPQBCqQWNFBUrq27W82cXzltycpTcpBpbG4PDXb5NT
N4EuGKY6XCk08gneJaUT34j72aum8UwC1mgFshFHtDjxkjgwQyPfWMfgp9EOEtxF
HozV2y3AhSJaCJLpjhoi1O754ij2D8LcgkFd4dMbIrnjFD1J5yFv61NvJqEzL4Lm
Sx00sgggHTxy5EKBQWTVagQOHnIYfviha41N8vQzo0R4NK0QS2jVviMbMW8IioJt
/yw71d4e3H0SMuqn7r0g3APutJ+QGGjSAZ9IDNHBXKZEq7bVO2kjbbVnmfapmS1F

`pragma protect end_protected
endmodule



module SB_DFFNS (Q, C, D, S);
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Lattice Semiconductor Corporation"
`pragma protect author_info="Lattice Semiconductor Corporation"
`pragma protect encrypt_agent="Radiant encrypt_hdl"
`pragma protect encrypt_agent_info="Radiant encrypt_hdl Version 1.0"

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP15_1"
`pragma protect key_method="rsa"
`pragma protect key_block
X/791CPQchd6RFFi2b6RnHuvpeuvdRJQnETHcdAMYCgiOnHJ0aEgtmNp8PzggISA
0554EWqa7O0qIqvo4iZV3XEZZPXiGt2+gbJ/fWbgc7bGI4byKCmXNRlQiV+wrUB7
FlrH2UhHezO9p3ArOr5sSFl+pV8HX7UQocSYLKVIONE7n6xJjkPbgPbaeNgUqfGC
1e0zz00WnvrwV+WZtRKUR5GafBxlbKeut+o5tMr3BFMyOmhmZCcIZT38qzuTPaha
p1Vl+tiUg8DcjsyBCGWSuDnvVtCcjogdSYESUG5ZO6nCOxYAgkxYGm7g364xNgJq
B5wfY+kuoN9ytHPKi++gYA==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
Mz3Okc05sRqziiF/EasEKBieyaBzDfYK/E00cJ3MhOBaHXpZ/z8NYAr0zS7rZBRi
xOoAdxYNRee7WYXEXuEPOwfWqLdKmH2KTNC3Bpi3l4eHgnfth8vYTo2XKuMnqOW1
vsB8LfZFz6DnHyz6uVWGl1XBRl9jQcHjZJGhwDu3f5mfD8Kbfif8HaC15MmvCJBV
JW0ds3kdNt6H+yhsneqDjqBSsXMS5LOzFA4Jg/Vp2GzkVA0ARTR+EBkaCnxSkgfw
grYfYVih+49EAoL7itn7XdlG2w+ef88N27EYp9XBmFU1PR4hAasRRS45+/AZGmFN
XIc1EXuw+duU3i0GNhO6xg==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-2"
`pragma protect key_method="rsa"
`pragma protect key_block
rOMWYhV2Ea5MWMV8MzqBQrTYWT5vL5Wa+wAVZ66ScX+6ViPj0wGV+5GxFnbqYFKK
EIvwNbKGg9/wBxKf3uWbUGxJIbshVJITsCs3r920R6sGk2bZb3N5MF4alb6jlDyU
yerKHiF8sJ+qFQsupN4f/DyZHSbaavH4ssn7GEgMZgVWfBDJ9FUtkpvauayZEjAL
/RQXUcOXeB2lKR0Ku6COC/VJ2XvkXlAC1y+L8zwaO3E0pG7uV/98+7gLpkNa6lu5
luX3YYEosy89W+yA7Rw2zVb/g+wkHSNCbVDWv9ZoUuLUvBwqJwhmNLFOccZ0yRmz
DhdmximxSWP8yrxF5PX4/A==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=128)
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect key_block
d/zn4hO4tWuox80mqRnXymZfAbX5dzPvlZcy0cD/3k0TS72d509VS0fK18dyh1yo
gTQ2Czajy29zRXp6gJ0WjpHz8X+CA4CxQCqyTXv2gjviB3182uXi6t9L0QEDx8ze
feCG3EEBDGDVdVsNQkiKebCyzS4lM1yeam8i1SCMqhE=

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Aldec"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect key_method="rsa"
`pragma protect key_block
VDUAsRojsLi2nukRtY09rCaPhtNoBq7JnB4+8Ow24U1tX9VNQrzO0p/Q6Nr66RFu
So3VvRkLeTJ6O/yTGToiBUWi0K1v9Qtatx5c/LIqhWf/fsHgUnHTm2WDBVwhzewd
ohZENk12USFSZXkWtV2BM52PrHNs9GhesOGQzOQi7avF+abl/CnCHJEwEUiVz766
R6IgljUe6u3BpyG3bCe3R+AnwTuX6NU16fU1oxViIr2P9WrOQuaRT/PYvXIFdIvr
KgVgUPVGQDCyLK/BS9x1ezbyoWUZz2YlChgE5I2rjSqXpHW9I1/O1EzSs2NdaHmw
BIAKxJpoxB6NtkPR/MSGGw==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect key_method="rsa"
`pragma protect key_block
hmV24Pcfnq9Xc8iQKmbLzvCDRfA9SCVe1PLk4l3iaSVEWI4FnoZJJFM4CacK3Bjb
LODMeErAu/NTrZq+ng55FZPAfubtDrmorNnWNbkreOUEopOhq6IsLzjAJiwb0I7X
h5mQIc1SdV7xXPYVPRHiVhvELxNhKrvusCqKMMupIdnsLqKqcLHZ+ILsGUn90dbw
oB88Qo6AGBxg1QZiIzRExTVLNTof9C6x5ULHOaONrkPd18YURcNj4NN2QiYTGQ/t
gYKErzuV7mBhVzbxAFwD211RMzxXqF5MoEyqfH+GumX581+jM6/7jSby43zuJP9L
kCEYlrdAKitr4/D55GK79w==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Lattice Semiconductor"
`pragma protect key_keyname="LSCC_RADIANT_1"
`pragma protect key_method="rsa"
`pragma protect key_block
XG2jeeRTP1HGi4E1UmhNJrJWr6vHHTdU4Y3wV2M57nJZFbO/E49B/F6x/Xxqg3Rt
/V6f/eu0vyoU0nBIyFBS2zml0YeiKASLWI5wkeBFWMbuLZxvZbsQ95Rli3o294CM
mwX+6PhxVyFUKpU6T/avxNHjdD16xeNHTL2iHF4dz+NQuWvaoaoJjPZrPWTtawYH
zCV4icJMnpZnPWPDFDC5WAt5CzQIsvVnkS8GiSAdN0b96C7GAc/Pm0pAokzCrqOs
g7GkbMu7pY8mHsW8+3eVutGdu67ipjtmPQfaUVh87hmF23stDSsp14h/kyAP+0jf
pjYiJNqoy109Rj+c5BS8Fg==

`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype="base64", line_length=64, bytes=240)
`pragma protect data_block
vTQpkpB1axfA1gXi3fGZHDzz03lhm/azLyp4mVDEKGd4iRDm8z2F6GZN5VD4LNHv
LVukO7p+9GVfIazsLhPBEAiMWsn7YrXEP7l6TQID3UYDCcEWFBksqC3Pku6eRPfl
i2qlfWodBkcoE3/53iC+4AvctsGzA1idTtsJmDY2XKTUD4hsEXCeHmxCURlfzf+d
hUTdIlKlWqQHakQ/NMXZA75vFXyQU8zhWxlyxP3HSbcGrWh96bL24eGtANFvmp1v
aOHdIXMLYaqicyqAAYNNh6Mu45++A3Ri7+sK88/Uul71xaLkPFdwuXYIhVkJHL0u

`pragma protect end_protected
endmodule



module SB_DFFN (Q, C, D);
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Lattice Semiconductor Corporation"
`pragma protect author_info="Lattice Semiconductor Corporation"
`pragma protect encrypt_agent="Radiant encrypt_hdl"
`pragma protect encrypt_agent_info="Radiant encrypt_hdl Version 1.0"

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP15_1"
`pragma protect key_method="rsa"
`pragma protect key_block
1Xf14+xGv9uackFRsgrchmo7fSgh7L4W9qJStdB+eUCZ7Mgia3ymGajsEd8OEi6Y
OVB76I59i7O76L5oWpLlPVvIov88F6Mc/kmO1RsY7R6wOdNQU5AC7jLjWN4R/djF
ganKPPKpo8lgpz+EdNRnA6N4wbMDUsdsYlV4xdEeM8wbXpr4eSd0JcJPzSLnIyL3
qceSqiSCLZmPOqV2pxtHU3E/r0/Ro2Utznkne1mMRCQ0+LxuKra/u4Dp5oNF266/
Tzrhk7VeD5lNB9NdGeCKz/cF1uuOKdcKfDhMsHXTMt25CVDB5fav9XIWNmcQZIQe
zBhqvKk1aPDH3Vheg3Y3rw==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
YxXvrBjXdqF3IjI9vaEyTK1zZTb7+obQSkWe6ephemfVYhC8yUkuh+c2N6LfWYrR
41SXgQeZUZeM5MXXTVZAbUiKLoFrtazhMLoxHq/bTf256EF9C4IaluGB50BA2Yus
77agDPAZSv3yo53QjiVN+C5tGs/OR/ElagnGoxqOrXDJc5QfRyU3C/txCrir5Tvd
QJnwc8y4qdVKDQNI3m6HBI12TatT1YAdXjE/ptsMWgu7NGJTp7Unwt706TiI6NE/
W86zS3flGYJ3vS1piyuAs0YOO0n0mbBXRYrZ0KyXXRaVZZ3c94OH/nqFq4ft1/tH
T4/P5WRlR96BfECWSLAxOQ==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-2"
`pragma protect key_method="rsa"
`pragma protect key_block
j2T5QAWnlcsXVdIfGFPm4dJ1OlzzMrN/3xCJ/i4t4xs+G7OFCQP6yw8uuO6dcMzd
m3eOvFR3cNGbrrMaD2p6IkQrGuuki0ZZMucuIuM/OxXDd+Hm9+jS4zHI+a3G7sN6
y0iotTJ37qLxFmbVO0uOqw8QOoowRdmKNcmcry/Bei2oI+TGTQ1LGK2cFkDup2gs
Ma6Ytdgqsk1nIVVeQLmPzdiXHgMW4rc8WIO6L6OfAiFDjmYmSfX84Rybz2ERfLHh
+qyqbxOAMOuVC8kftD1wk+kqn5V2uFn+aj6QcvvFrvQ/+hXxwuRQPdvybFUebnKD
q75IizSJ+jyw/q3O6w0xcA==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=128)
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect key_block
kWLuaQIjGldLmC7IZu3caLy1dqhdZbaHUMo8kCtipAjD/0AAVWI+1WyLbDJvkdJK
rpJwON860CxDuOUlkbsHl1o1BbYksEsMaT7uBArxvNeMlntneIT84LzzsZyiUUdR
tWUpU244jr2zHWcZDtrH7no6dYq18WkgtY6QRlCJg2I=

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Aldec"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect key_method="rsa"
`pragma protect key_block
a/ewRMRdUx0GdgXdE7HmFNFMpAmsUb7GdIdoCYWN0xczCSPJQZZdn+++gPNGfkTK
RLWFYIG4OWoGlyeZgjc6aghCI1Z2+5oCQxcSpsnNOAWIZf2J4NFnOrFBCLF/A7Rw
rcO8LMSqpLdfoyI5GpdLYtiW+g+kl67/hIalAMZtKWYheiGVxmthYqLG7QZLPkjK
98eXRFGm5WOlU7+VB+nfauUhhAUhWaVxEqB3ACRQFl6lgiooiotr+xT8Tb0HmEJP
gz+KEKd6HalARZS8IXPAMH+4vS/RpQ0XnUnhlvFJpNyIWeIGBe6HvD6QdQ2wsyru
xmotRYjn2hwsLPa5XN9wYw==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect key_method="rsa"
`pragma protect key_block
jJW9o3Xf0/uWjc2U0ybcagAGlnOGv2lwAmfEXE20Xd3wFdaS5WQrhgDM1zursYfq
TL6rcgyvPl1D2BNHLf8YT3Rhy04iRzNNlqT68kaBLpS54X6YslmokbaFZ2S9sa5B
reOWldT1SnaStxqjGFwoEIQykURVxItrAdzdqW6XBZwu9IwEA97ljJLx7kwl/Mu2
0/8pFD418C3cFVgooKyNHZK6IUCzihneIRmX8B4wLwKylAr+dCOw7M6YHfdvr+81
3B8UhL3FO0jUGxSPYmSjHQIheCqmPadUdDXIjzDvKfEjbYdk+lMVQj0grdZA+tOz
kj4GC4nktLSNATZJZhKx9g==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Lattice Semiconductor"
`pragma protect key_keyname="LSCC_RADIANT_1"
`pragma protect key_method="rsa"
`pragma protect key_block
jyEwg1fXx3cUX7Y0biuvZCnsJk2GJmd5KxtMRyepv/1xd2EKq8j0XtYM/Hb3qp4Y
0ecm5X0sCEzM7Crt70L7zQO1ZvAfchMlJUHpYIHXbHh2PbgPqeSuu2/tshX1NovF
8hHiNsI9KOnJSh8kz7+739Zgwz9iI7W/VUMAXOrabSXaGHNoYL2MUBAKiFmuD56u
UOOi1WAmxGpdq7dgAlPFBUjylNVEYJv5UHyvnJ46/O35A6uf520BrMDRxV0fbUro
VabxWnjO4I3mHQ/v9JESHqCsqhYIuyuiDenwXXfI7FipEyAe5IfaFkbEuG4CUfXl
9I9XZXhOfw2Rl5qP6RAo3w==

`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype="base64", line_length=64, bytes=272)
`pragma protect data_block
1+79e+dCyHfHDk6Mjw//oMqdilL9J08cQgOVAM4MWy2G9LI62Es6rD8cE7cdrT5w
9n5bcNTK6nTMbmfjqH4dgZVYFdPd2fzeDKN0A0MHJ+i/FQLi9utWu0viFhxYJMjQ
eEG305sytdqhj74S5NYxinPJDD3lrDjIJBvas77yNUHFtgxjVFINviQsi7Yyn7t4
CCYPofqksGR1wQ/j/AdFmpj+r0tia6E/3TsDQnb+0pkR8w/caS0ZoEPXyoZQsrAg
pjd5lEw73L+iwZHhEGAhZVLQ4nVzs9PcMuJWGsorfNWG586+YY1ke+9mqsz4QOmz
93TmO/RcPQQNArxsR1zzIhlYzjydOuIsZSTubKLb+UE=

`pragma protect end_protected
endmodule



module SB_DFFR (Q, C, D, R);
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Lattice Semiconductor Corporation"
`pragma protect author_info="Lattice Semiconductor Corporation"
`pragma protect encrypt_agent="Radiant encrypt_hdl"
`pragma protect encrypt_agent_info="Radiant encrypt_hdl Version 1.0"

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP15_1"
`pragma protect key_method="rsa"
`pragma protect key_block
CEi5ELLMgDma+71tVCCMDrgOejqiD6q+6FNy1JFCm0jfXreEwZMWOAz0B29DUTxe
mF932RPLouzX9wkMF8xJNOPf/J01XVQ2DvNAtUSM+nrmRTUPA8AYVT4B24sU5Hd1
io7iK9OfBHFGVlUdH34V4ncajUendl1TnnTTQ8otiNSB26vFde1pCCl62KcOnu9V
OuDkOCd8tm6au3fiqnZCllfEN+ehJqb4t0rGN5Z7EfUBNffQcgMC6RF8qeug3pOC
plXjHbZSEAseNUWR52jx2bmPq7WG+R1bjkO2PEfsAZdKbPZr7xUP0kGI7rkSrHhW
CARBzLwQbsPUn4qiNXl1/Q==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
JhTGSEnKhePORF9e+WCF6OZxxCH6SRArNB5h57gO7+21PkSKiDtwF2cGPcIL6PUa
YKAvuaxv+S2MQdOAQlE2K2gnh/AOrKygc7Vup4vNUsdpjvF78e6IUwAUsBwgNTAt
vlWmqI+sknVaQxZ6xWZ+hkr/ilFjeiQgDJh6lpUiEzuPxm1EqTQqjHksxJcouLqF
t+yT/SYDFt/ep1MINHVB6E1tOhTXD7mmTignytweVqBJlT8FimDAUHiU83+rGCoo
YixgJa5zDRZNTmYk6dDnMp07ZmEY/fsbRUD8bwKnym9F2BL0V9VHnw9Z1sqgYgyW
/muPAp3CEzhQUBtw4lyuFA==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-2"
`pragma protect key_method="rsa"
`pragma protect key_block
kYtJSvATmK53pyD8+CfS66R02HtqEk1ONcwpfoG1qI7eD6/YR/5pSL5IwrsA444J
B9wA8fd9AJl1gXSQrsPzCV/zkniISOCz9U/5mY49uJXaUwjRCCD1V/u+zjUAxpI6
SDxpCxTfQnEJR+lReBT3vqTibjnP04uBFGapimmti8MArjqs9giM+tYw6T+YKVv7
w51GvMZhqFHRG4ckydu6BydW3BsIwEVXfyUTJ4AQJ5gKrQpJjkSnMS7yFC/Indb7
0v+6dw77PmtoJqjkL8X38YYSmyGRKtSTl9oDVgYstWOYIB5cSPQveM8ANA9h8br2
Pk5Bu8ABEeDTIBBkWhp0eA==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=128)
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect key_block
RPfvvT8efQ9+VrZIx8uznNfJhvj1T2zeyXrC5ZcQRGOyNBrAyKePmR/CyyaEZtAb
2EQOh/bTfEYatlgsHMapC5biwxo3wnx64gdl81jc4cVM56aTWZdtAgvRHAfubzCx
b82WBbLn8q/+fZdwmzk6HUMXeQGS6dbu/5tZRYvsNG4=

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Aldec"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect key_method="rsa"
`pragma protect key_block
aJXzpUgpyg6dPS41LXuB3DrN/cOGNuokUtoXGHnoECDhR8rxe/ur+RnwNdAQ7RZr
YJnH8On8P8J/KEY7UFEvmM5itcYigsqS7n4qQ/ojRa+u6qXR6K0fD/ywMv6KihYB
/TD8oIPOtFtEs8eLGx5ExVchUA39n2VPaWDf004a1GJUldHLldb/XwBPiloSHzwK
SPob50AH3ECs74UainqYGpqypHyDPNUOh8Whzj5K+3aZNmqEdGLRLzkWKcXP/zIj
zJi/yB9EpX7aDmxgvWcMo/B3z11RWgrH3qpNii0q1a7wcwG0JmY2ENs5FMFxjLIe
dHfv0v8mTpZOqkc+rpdXpg==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect key_method="rsa"
`pragma protect key_block
Tg4NAwz6BD0kw3JtUAlAynHgCw+R38FhXxiBo4yrLmPVTjDAs29z+DrW0cbPNgy8
nmXs5JpF7z+GlphR6vi6AHaxMAbFDHcHzIJ8GHne16Sw2OiORtxy+S/ptnOIXALu
1G2xQS2BUj+w5ZdxSMUR4703tDkCqdS+n15FPX16ivnNXa/7WJdT3z1KXb7hMLUF
VZh+eeJmonimPvCba1V1w1Dl8UrhGbeE7Eug74Kb0vvWzQKd3GuFp4Qz3ibSxxj/
2YlyqM0m1YuOoCAQqP8sofxi18ObZmp3mrbiZXHt82dVYuUHsSnotoJr2AmjFNgD
/EKQTmg8mCASHXzeipLwfA==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Lattice Semiconductor"
`pragma protect key_keyname="LSCC_RADIANT_1"
`pragma protect key_method="rsa"
`pragma protect key_block
DQApA3rsFNxulnIPiShkLKnQwpma2ACBw0R3sDjtxtAuGBxMdaqcW3j/5UU1tUdj
vXJufChcgYaj5PsqkFh4I+CP1sslv2ALsfHhi95db1VOVP+Tmx65DOWy4yNIICjp
F2yxddXVVym177D/RFRXR3BLqEmBt/zi6c+Qp0eGz5YTfoOmh9dFte9MRzLdZ3xM
VfF3/WB01Of3LsWIQWjQ45SNw9lFJZhQXp0KakM0IDavg4HBDexTCII0XiIvmvt2
oHv07FzTy8eS3ck5wqVJWnUhJLMTzsjiHOkuaSV3hOS3GfHXJWd0/8XVzjL0PWBv
DLDSs9F2IFXMkkqNVa3qmw==

`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype="base64", line_length=64, bytes=208)
`pragma protect data_block
zutzBvCkSYI7a6uo49c/I2irBDubl7k7uDrg3R+FAbzU6MWMamx7LLfzUnhZLzV7
w8JxaFbSDLOdb6PFzQ7HknE9+xUGrNTvNPq0vqK06auvHtUtsytCROTXF3goS0qy
z0a44juk7t30H+1P3zmgCrYYuCTqO9UBO8Qe3n7+7Y3b0c3QQyM2rg16YvEMmiXx
WKXmajTb4GdwUvoKNxnm0ZOFiYe4hSRCBYnP0QKe+jcQeWl6eu5kwobM3MyaLUSU
jc0HT03Jjh+27SSfCZxGAA==

`pragma protect end_protected
endmodule



module SB_DFFSR (Q, C, D, R);
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Lattice Semiconductor Corporation"
`pragma protect author_info="Lattice Semiconductor Corporation"
`pragma protect encrypt_agent="Radiant encrypt_hdl"
`pragma protect encrypt_agent_info="Radiant encrypt_hdl Version 1.0"

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP15_1"
`pragma protect key_method="rsa"
`pragma protect key_block
Odl/tykRG0mHiB1VPeIAToa/x7cnthOg1HvqxDXwkkWCCHOyf/QKnxmNcg1hehbl
PvQqYkLDWeVvbCDFd9/qpCYgHvIpYrz21nCfIhr6fZb7RITT1v+II8Bd14qefgyu
mngCw9fdkmXFx5+mE1TrGtV2R8hdZC3kUlBMszjFPcWZxVOhM6aPeBrxN5MojhnI
yu321qhzMD0poCigFw2FnW0V8d0GNYaYpTqu6TGa2XBbxw1n8PGQ+njqL/A318Js
QZH6xsvThICGWSWs7U1vg7abJcCjp3kDBVU2Rog+tnOFJ2CTd8zz7uW1TCG2eucs
jCZjI6bkldsKbTRb3aAzdQ==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
VeblCHZz+EO+WAK28vZHCrK7OnTIxR9ldEcUciAG+jykdnbsK/rxcvOhsdaqH6Ti
GoFngJg8v1dXLWnTON7DfM1z4w8yKwb+t+H6aAGj5O5lmT6DF2D3JcMJMofUSXQj
tlENweWRdA89tjDWqGtvFr3PRYFvqaX3YPg01QBi0oWoN67jKbIuFe5s3iuaKi++
APcoKVM9WxqsByP6QkBc9jja02yynmtUK0RQ4WP+aE70yNlEAtZGgA35R2V5EDLH
8UaNlSAKrf6N8qGmNgTj7RftlYUYQL815D/ati/BvlHDClKu2fvxenZD7FYvMPOQ
QCHO5Dtw48xgFfUzGT4Tgg==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-2"
`pragma protect key_method="rsa"
`pragma protect key_block
SG2004gZ7B1mjF+SXU6PpJkqA5bsvqlYx6+e9O0EA+2FccYZPhvcqXk3vO+LH+HH
ASqrEoXaatm5Fu6+OPmcQTzVNhxaFMb8iKeRlqWrxMhuWxshIsq68xG0lOa66C+S
w71JyrQyDusa+fRQ4HllOLJd+sNl9KE71B/qCFyYxR1qOSXVkak/CY/w1CrOxvz6
F9YRrM+RJkusRxhYK5KfIavFMtvCx0dtwT0BTHiDP6LUBWBV1S76lhI63/2T8W7U
SaPm2+xZuAR2xfXm0Z5xdVJim+p5b6BKekjnHFQyoBvQJJII0w/sewJKUO6y2LvM
s0lIoTBiMQ5J54wlqpz7cw==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=128)
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect key_block
kMoqXvnipsV42ZHTAj1ft7jXZfu/4FCIURCjnf0y10x92/J0yjtbx/dfxMe0bqRc
qwagJTMFC3gm5yBGAe4C9J56BoHmZXLT5HhMU4JTwKFney2o2fuXhdjg38H7oCUb
xUYij93vB+NZ3WLAPL9GMiYxR39yLKrs1yaWXOGlNRw=

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Aldec"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect key_method="rsa"
`pragma protect key_block
f/83yAwmJTGuhk0bqG+8/ll4rlzFoBp9HTd0sS2L2bAXZBPxywB1LJygwtip3/WL
m3qMOwHGFV31YEEs9GzFRpy5Hvivb6mewdBmB0fHtstW6KksY6YnuzdAHN0W+4DY
0d9OnLtBbaRGQ5NLYlu46QkkNsF6BcRuuDfQYwIg7+T0nxyhQCJx1+e6iwj8nfId
z49fr3QUY+i6SjYezJhQiR56ADjFjSCWQnBUZE+NB5y6ZGnveCjf2/3ra74WGH5k
W9ZCqssT4U4hAye5/YDkYNpyPpw02aMIp6mjwR8TWqXf5zgO+B2It0i1zxJ5rHrV
Cvvd4POLCLg9p3tZdbZkrg==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect key_method="rsa"
`pragma protect key_block
ZhnWtedkg7Jh29XCRYqyoytrKK52xA+xfmOTrie1SIn/FKULSiqohQZ/EoAcX86C
vBK3ffvDeDvOrqUL7LjaUln5H8jx1KXc8qumyHELgwPdRpFIxrdFpCwJKG59gCxB
SYcrO1VMHe/WsqZ0dII20TUGT3qu9V8nHYOyt1JO8RmwIz35hrxnhd2oI3dEn5nD
rRz0eR7QPBGauhh1IBMaq87JDweaZvFUmZ984CM9eEXyv8KmKTk4H/3gbPEaxI94
BQqbJFx85hycvnZoOPgGFfMyOeW8UXPzGFznVxJHDFL2a/QaaHeH4VXJdtewhHuU
LPNeQI5k5sT6uZG7rPacyw==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Lattice Semiconductor"
`pragma protect key_keyname="LSCC_RADIANT_1"
`pragma protect key_method="rsa"
`pragma protect key_block
le+NVXunOe6HWlIGXWE4FgIJLAxgGcQL92afgwlyLHepzCCuMDAfKs13+0U5H8jp
02D+fBDwLcIqMP9aSJAvmFuRfXtrZR9+/WrJoCA3DuZzLbYVtf5UOLc716ithJPa
m674/K5Xba8Jf5N2/hKFrZ4GW4vqAwXXvro1N9CMHx6/a/IH6O1gNHdbQIchd+uM
2YvSzDgjyYLHi6kY8PtzagKa7yKsDs51BNFH/z98ayUcZSeavqbtW0XxfQjL18qR
czhNf0WCGNpw5VAOC2IAgZMNhIHkBI/1T35tNQ174PmMGtbA9fLdCja1PJG6CnIN
EHAm7b+f90l5d0offHhF5A==

`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype="base64", line_length=64, bytes=208)
`pragma protect data_block
iG34oj5sw/klgPU40RJeAAgKp+/9INahyfdaeb+jFoX3bJ98MY+352kPWLgjLMOp
7oDWWwQwhYoq4tofiQIDlNM/AwSndtpZiOA5c1tza/k3w3AasnXGddjO6wkG6rhD
OAfY9XLgnuzrZZFcE3X6xbscy9aEhS6Ho6y8Xjus9T/LMp6WmKtmDS3t/DK33bOI
I14CiiKhNk6XU/lpuRUCVD6D8M5wyUeaN3QWd/15/lRcotov0Pt++RL/OFHO2ko9
GVtd73UfQI6RP4Mpzm+aJw==

`pragma protect end_protected
endmodule



module SB_DFFSS (Q, C, D, S);
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Lattice Semiconductor Corporation"
`pragma protect author_info="Lattice Semiconductor Corporation"
`pragma protect encrypt_agent="Radiant encrypt_hdl"
`pragma protect encrypt_agent_info="Radiant encrypt_hdl Version 1.0"

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP15_1"
`pragma protect key_method="rsa"
`pragma protect key_block
1tGXbZa1M8JIAuqK1PybK6TLNxe9dtjjbdK/gOIJZVy2d5YuBVQ2215bxXJHqF1i
deCp6HoWZLjMr4xcZSh5BU1QoXVuCeQr/LLlOrU014uIbFlboU8bJJQ4ay4PUje2
8oXYzq9TMbu7/4K8OcSOfo0DrfcBieiHkoNiutr4dwDYPtRMqF2S5TJa2Byu2Er/
zUzkhGCvSU1fnan+3Y7vKG6M/YKODnH/jWwfuojmsCgkogEEyx5g8d58+E7xSRfq
PuScl8/V4uxWOcSHLwkHHz1njbCaJhGB0cRhBSFQkCf7rRcz6s16F2AdH0G4vKam
zU5UDOFfcFCABWFoGCEtIA==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
DFMUAy4/bEgIaD5693y+e89jOKsyAQbOwN3vWKG5lxlaHsGnvsO4pt1Dfl2rlj2K
V69zkzcUUdQisWCWCplW6rhVqYowKgej31ctZYJDkc3qxErIY7KMqtXdT0XqAXYd
ql6OiyUNIjbCI9AgY4sGibAQ7birTK6KHxK0XhdPyN4xm72jiIsV/F7/6E0omgkl
RQJE+D6s9qUP4O1Irt28OyQtN5381/ngMEzwBCBmFv4WnVJ1Yuie+nmulMkkdExC
GOW+Q1os9ilreZo+HGnNK1H+1sd9xH88SbQTKvw3B+j7hJQWwveXl+hEoIpre4zI
2kQa11UaONX7fV5gkT9CRQ==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-2"
`pragma protect key_method="rsa"
`pragma protect key_block
f3hEPOT/h69D3mJ/BFjV4qo+5zkeF3JKCMzZS1YTsOfa6Sc279buxUxjoV3AAHzN
HKgK9BgngFjIqCt0Wfx48MZQR1iOMq9Ptsxf+2pATzLIkPAad5sF5yUjgtqmkyfs
3Qqa8YP+jsbcHxfDWRhR1lthuEZYZRdMd93J0Kk7I2pjhPZBHAM+jXHIqqojicEh
3hjahRQLKsc/mrVdNdqVhlpjozDr7iGD7bVwcSspLTLGvhlYmJ5m7/Ue/h+5OI4u
J5IUpM709nxgdpGZcbxN1bLCIMVe7kF9C2NY5NJ3SeM+ev1L3cMsAClzr9sJy/0t
AF597o6JVcx40SFUSymUYA==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=128)
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect key_block
1b80Qm8j6Ukx8w9cGDFMeetcmBl8vW3DkQL0l3HD1Dhw0gorIAv0o+epzR7tszto
dz+qiEh+Y9/K3AVoIqELwg2tASz6lyDAuNyGG6FVSCBKIU32m7fW8MMVECBAy32e
acaMSGDHWOHbHwyAoLXo13Zz9VyPyUVIl5tvD5bTNcg=

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Aldec"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect key_method="rsa"
`pragma protect key_block
lpLePOV327ZkrLzjBwd+MGGUMHoyPHzZGKTdMHnErii7R4Ep0emEbNPZ66D7cASa
VMQCkcyyZ8hnc8lLOGl6XS5RUe6gGovXOD8BUQQeDSILnVEm4V7L5gQKnbPB2xig
1R0IO9ycOlgSnmrVblEI54eUzOzAGX6eOzCiFqhtFl1cJxtUrs9T/dSWvN+gmIDZ
Dytym39xwNEmKRqbdYGpi9Oj2VH0WY22xG+YLfE+ENQYUD4/wSsuxnaS/Mb5iHfH
qPis8q6cp9/L6pYHlAYPvZ2QcsPH3Xs1Z3w1aUvfqHzTpAv0J47/411OHs3eVwQ5
77rfWEFqEAyLWPejwwi53w==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect key_method="rsa"
`pragma protect key_block
eEwRAm/zkSIB5qI4o1SB3vCl7ZJwTbrBAyNI7/lKHOJYSDIb7Q3Q2e1PrCJwk5jf
JmTdrqMmUGFSvM+5tGTGN4eR0PttUQRKPARG0cTTnv3onfcFxmpBx9Oxo8TKkYWx
ei0BllkiLxpCkFFTZOpGj6SL3gVm8NmUxVb5ySBKcpyw2yllM3yZhKIYbP0XTmrU
ZuZtcwi0Rj3LI656EdbDzi7XrxK0cGHN5FfoiwoYCR2ii9knNMzGh/UHQvCSSbCL
lpaH1yxltT4K/h/Pqu2mcXT31fewS+lcP/ar+q6ahMUwJt/0rEdEbhNRDBTeNlEa
C8cLzJDaTtIDAleBnqZmzA==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Lattice Semiconductor"
`pragma protect key_keyname="LSCC_RADIANT_1"
`pragma protect key_method="rsa"
`pragma protect key_block
Z3UbrZpEBL48oVkEiSz3enOuxzq7Pu29HjGvhuiW/1f9u0DhWVTWbzTAUaUzzjyS
zdDTH5Cji06hDwxaS4ICeGYweJkbUj2Ph2C9O54o30rwsRSYDLukk/F6/3G4ckjB
wdrXsfcuWNC1S5l9CixZY8Cs/sj3f9Hvw/bFeyNLVLii8DQjWB6s71tqA6GHGiyb
W0SEVJxfS8b5FxU34qx5uXxO2BQ+YYsJ7Pvp7GhCWeCXH9AsE0bmmoR6w+ayWlth
7ReQJNUyG69zNTWFFn/pRtRBCj9edkkS9QH6Xo2+G0JbQYDhOQJkAlcwTNOs0dZv
n3QdEhe8MaiI6h6W2kLDWw==

`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype="base64", line_length=64, bytes=208)
`pragma protect data_block
UWmt+nKMZbhmlfKTtnMdvIdy8Ak5HxcirOxOvtrwEgD4POcqjKDm75Ds+5jkGs48
c026vEPjOxEOICE0TYrb7yYwk3DmZZjFT7QTzex9QXcy4zdSb5jHVaTF+qiJrmoW
nWHIptGQiMOZULMAgsLl9grm0xBPTzvGbwt+JHoh6VqYzyUTICiV+MZjKPx3rfre
PKriK8q8AGi46q5eZ1EGgos9Sikfq3uyXXRZNZg4DME9DibsUBeAxTvXIxQamedy
gG4Y3hfSEyZGDxaJUdCXNA==

`pragma protect end_protected
endmodule



module SB_DFFS (Q, C, D, S);
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Lattice Semiconductor Corporation"
`pragma protect author_info="Lattice Semiconductor Corporation"
`pragma protect encrypt_agent="Radiant encrypt_hdl"
`pragma protect encrypt_agent_info="Radiant encrypt_hdl Version 1.0"

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP15_1"
`pragma protect key_method="rsa"
`pragma protect key_block
KVQ/RHbrJocHFagcQEn8vj2YMwXomnK5EPUjd5E9cUAhh0sWAD1uMWNhXW/ElpVW
y9ZcxRbJDnFjLTG+2T6co4TYRHhjsH2RyrVTvBTvGewkLzwFWwqUiY7JupQdaUcC
YQ/knDxsn+IvTcWL0wL8oe9DwAvEUuCQtwzyFHVMW56soTomunU+Jo+lTI2eGyJ9
18yjlvoCDMD4yAFE10ymsnII8uppPwMxkEwwf2s02vx6A7z+L56yJddQZ+dpp3d8
/LBopWLlYFSiqvXF0Jt7bURuX21T5gzGBywSq0B0vxOOlgPpP0fVKw+Iso6b6APw
e7SFWFDL9ryiS6LE4uK5VQ==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
m8NMfI6/eLX/zSAiXshn6D8Mx5XYpxc7pCO9ZVoBbvugoXNwYL+EjhvoX2801piY
Ldj4q92l/9vX6tNsuipHamuX9ESGOoAqR3PXXb/6VTaQWT2FezNVORS7osvCKLZc
to7B4ERe0WBE8IgpJ3EomMBIh3VyvdKRHlRk4xKU2I5kYOvOioK7t7bZjj3YOW7L
jrpkPfx7t5f+GHvICeHlh3DWzKsqK7KO3OUkM6FSXsc6yWCMvGC/HagaJPbB5BYw
wc2gb29mMqVw2YvWNvk8I/G15lfLcc9H9MRb0QRgrQpSh4Cu5vD92RB4q26DpGbS
mm2lB4QWy38/E3RMex8QZA==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-2"
`pragma protect key_method="rsa"
`pragma protect key_block
noRtjNPHIQxzP/LS4EWZpZknAVkVZZyFECzPnorT8OY0rUtSzapP1l18bvQTWEQV
IyRiNARpqgnVC25dKt0phbk/hZUylSv59oBPFdA+Ls5qZuVTtmjO6vgN/yC0p0wY
Qnqz+royMhSPQvcdAc2CK5YA/oTAs08s4fJiYcnpdsW/61Jg1e42c7U4hOmCcREp
dPuXXZ465AzjwWIe2p5h5m/NzhNIAXM7dIn00wy8rIuJGYJfBaEdct+He9zIZkSP
bt0K9LSiCwsafXemqZuXvq3eSifH+SiXav9/v6v2XuiA7EFB++FwP/XqpJOmQXTQ
RDnQJOvnfCbRqfMjtT8Zbw==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=128)
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect key_block
N/YBV3XM1fJA2xeK+XTVyhgJHB0+U4ba465SxgAytNVq9YMFiM1Kph3ukEJztH2P
+6l2C4kjv6zf4EfCKsJKZMSDPdYnNOD3RFnTSxo+C4//11GextgId+atXKAaUij/
O4kcI0goZn5tigMBFtexxkQsujpz4LrQlhO3FJ1zS9c=

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Aldec"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect key_method="rsa"
`pragma protect key_block
ULeyqwqwGtVhNIu44dZJXT57cNgh8Z64MiECc/rWe4+2zBm+tW1GY1OAVLglIbJ0
7AdCclckdaQJfOO4zbYQN4VieJFqZm2tZ7ruoDg3iCH6vW41l0KnEjYD9Aherrwa
+3eZBDEDujOQlNl2puy3pXPNNuBMncHjvgxIbj7O5KayjrOMYSaZf9Q+UlADlIQ4
UzhdFX0eJVFG8tCuMDFhMHCLAWCUl8u5PipdM45rthKd1cMmy6b1jRY3I4/JyGqk
Nv1mPyGGKB1ju30ANDNDKc/M4GaO3X+2rQUvGpO93X7ldCYLbwxJK5JkLJ1ymRQ2
vojYHCJPOMi5QOn8DRmSrg==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect key_method="rsa"
`pragma protect key_block
H69+GXOFGqjS4TYKDs5lJ1chnEI4a3cjRZqjQ+t8+9usfK/paPMC55qLmUfZjU+w
8McEb44jO8csLlw7LRf2qZuCGLScEJw3+bPOQa+HhI1Y8dK38CDqAcBPiykdZ3X1
elGZ9w9P4Gq3YqDyOtgpRg57OnE/fXj8TRt3FvfXEBkCI9LY3pdkmYQqrpAiIoBn
XggFbtYjNaUkvvnkfl05sZxUEOM4Ju70FMMDT5taXmWKMXBIB9UOJKhNMmschuqO
vh/KiScZPMxttxnFiIRZiYH0wN+xjA/bVHbPxti434okVXd+4cem7ilXHaQMweKp
45fGomMKkY7dkqS1x4wXfA==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Lattice Semiconductor"
`pragma protect key_keyname="LSCC_RADIANT_1"
`pragma protect key_method="rsa"
`pragma protect key_block
cvzEcJj6dc6HzhAjd1zxEjbeZDtOg71G1C0DqR4SS2b6El6tUxgmNFHbMTIiG45m
swKZznp3SpAG9DdPbGdQU7Ja834a1As/8AMYG/Mx2IBYe+kjJR2chVozSlBZQPQy
hr0KcXblooAltQ5MSKxbXQDljnILHKfaOzZHbCirntjT0/+6OEAV5Mrqs3789MXL
JJ0JiszPYTGrAFXoRHgqSktJRaqv/qKqaHmBFCd4l7YT1EEs45/HvIdzuRz73LbK
CnUkHEbLcDcXd4iHc12B/tKCdisMa1QJQgSBATGOOp4kdJN5yFMlCmvcktj2kXYF
xRbwXB+N15OaHx0qNSuPWA==

`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype="base64", line_length=64, bytes=208)
`pragma protect data_block
wbN257RcDFrzMojpAmoje9tw6JN3YaOIK6ySLvYp1SqPv6031wGGlATBUEziTkf4
6+SytVrY0xHfLJS+wrgS6Fe+RKge05tMe8YpkFLd8r9ere0vBuEtW505NI6igu3r
qGhN+LJ6+sVnANipGwha9Brxq1FNDm7gR4fu6Fs1HIsAJ4TLuFrhaUiWUXX+nrlA
imijmkKkurZO2bC+TXpE0Fs0ewqUrpTbCpaXzsvuGlonykkZGt6c4lWqSrk2+9BK
nYzSe+LMSSVmaUdgfUgroQ==

`pragma protect end_protected
endmodule



module SB_DFF (Q, C, D);
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Lattice Semiconductor Corporation"
`pragma protect author_info="Lattice Semiconductor Corporation"
`pragma protect encrypt_agent="Radiant encrypt_hdl"
`pragma protect encrypt_agent_info="Radiant encrypt_hdl Version 1.0"

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP15_1"
`pragma protect key_method="rsa"
`pragma protect key_block
Cbc+KhfTg9tVE5UAaU2k+MGegZwF8ynwN/2ahyYbArHo3sRBDEidEOCTAcKMZgMD
s4tbcpKX9kOihQOOsS7MKR/PQQfjb39L7f0SyXmqflOGhsMfeOy8wuAriq+OJKf1
uunPsOk6/W6lhPvEL3/r762pEnf32giHvZd1JzemJFtwUSVvBAtLqWfIG7WGt7ZD
F6ZjO5ds9KtwvV6Zbtcit5QAgMcmBSV+LsuM4GZxMp+P8Xz7GiYh8xnSnTb26O5t
DDNPhWE+HwhNszn5rcMzV3HisHI6wgh73+gDHqZfKtMv7dRW+XRw3UKR/AHFML/M
GjcywJRB3wqtFSThdOMTEw==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
WGg2cnox6YHJVov53MxMbANUL17VFIZ4D+Jm0OJ7dsPeeNk+a9QBWz/gaBiKAfPj
gN7zxWUwUNQCc5uDj50m/wQ3k2sfHD+vYIw+CNMsDnRarWrMCBS1JJxNWbOlAOwA
q7Fx9PzvM4u55fsi3Ld27gGhDU29sYbtcMNTgq2L5wRxjQ+WLddybn/foTaYx6tX
a0PQ2IuOABWOU7mlXCs4zEjYX48qLSCFsWq46B6rFaUbZb5RHSUqlNxhKOO43SEE
heng7ehT1BScbyAVkHJnJtF1oOrDLRKjLh6yhE+AjP+J+H02UGgWAgpB3FYnaPsZ
mcnUxnsBFnzpVaCyO9Hy3g==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-2"
`pragma protect key_method="rsa"
`pragma protect key_block
bY+Hh9Dj4nkCCDIgBQpYRucWoKi7JD8Dmx9REtQWfThX/b/d6wEGADuaGq7r93FT
9IwfQm7Ie/ktk49Zp8LL7CIlRmFTkeJZRtEyVFTERQ96DCzh7QvunvUZoAymQ3Sr
06CFoKG4ltROeSfy/wDxB8gWG8500fbYhmRKFIM2UlzgGezgAZEtgQocxkqAOjoH
Q1YFnIHTni9QmCdVfKl1RVbCDPeTj0Sgv/Y9Tika6h/2pvnopOZF1wMNfvIF18ZA
SskkTbjqreVPz54JhM92bCSZMv8W0G2nWsYlcuWDegwxV2vAGg0jF0HgADm2o51j
IBaIMnJ286+CdgpHpI93Gg==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=128)
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect key_block
QJLxe77A+8z8+cd+12opJ8YalbL5qm8UYgoDeu5e6gckMgpw3qjYNJjaen4hRf9x
LfsW0zrBgJUN4PykahgFLTlrqt9medt7j2UzLBpFBOzde5jevdwZCJEMqte7eN9p
oWPs5R2oFkJzBfNf8i4qGfawqOUWHLR0b1LKTNEYrJM=

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Aldec"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect key_method="rsa"
`pragma protect key_block
kGKJYAoBGMSudR+V2Kyk9fwFXzzr6Nm66+3ajQDFZnOzTmZG3uDdvP+WNbmD8jPU
FumUQcreJVShTkJPQnhoY5rQHEi8y/ngfRp8kWraWRaE3Xv9X8ewru5jz9YvJ5/q
0txd6PYhYtdH4U3EsQvv11BxJ7sSUX0GZ1zFd2Y5C79HJ3he+PcZM/8f5nkwMeG2
fXNkUtJk3ZxkFTYuGcfzX795oD1tt4EBNbytT3b6uj1kcPUdu4H/xT08uaS17Gw3
xqjF5NHzZkY3VGaYW9PxIWmT6jWM0FXCYV/QqHhivoFlFO8BSsZoWBfIcb2Hz4BM
E9VDQ8Cz/DNGrEsFOIZ9KQ==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect key_method="rsa"
`pragma protect key_block
QVh+P1ZaaUhAfD6Hb/v3akoRYaWMJZJ7SIrtQda/FlOOZOZ8rHuBc/aF8JzokQwJ
5RZsgfN+b7RepBRXvxpA40aKVCitCKXFCrkmVXweERrjai8d6IAevAOBh9nJn0Se
mmUGQ47X0HAWFm4vq+w6rdNzS0QvECu4AiZZ33jfDQGJQu5HeVnQo45vx8W48ysp
trY94m6EEm2m9a5hCu5PmU3NSmHKCrUoaL7DgqHPYFYa1UEyQFh+ZJNMny5EE0dB
bgU6DWV4Ho8UNadPd3DgcRYp6lS3Ux6xm+Q0UFqr5FN5ItWZcE3XlTNHKzBVfLan
LA5HtFbbzQFX7jnJj7/GZA==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Lattice Semiconductor"
`pragma protect key_keyname="LSCC_RADIANT_1"
`pragma protect key_method="rsa"
`pragma protect key_block
EWpX/Gxf1OEqaQFBiZcGUaN8k2qc29lpmL2pE00mfdPxuFDjH2n8J/3y1HgX6T9W
fsk3cUhrDCwBPY0OGDAoD5C7KKzrvyWt0INUeOZaii8hA4DmLAYaf17S3Drtphja
efVX+Fx1IrmqgqtZ4Tjx/MTbXckgrk8u1RM8vSAzeZI0lgJSymreOvedOjD4rDnh
Og9by1TSa74Muvoer6wxzYLd+8NFE6xeEUJDuoU0SRNt5RmkLTfLvXLoYTVwVIue
ZQbJFIMqCuoqvSWMS3ZaRjrXFXsm1GCm3pcloNjczOcc93cq/YhR7zMxwbOBu1mT
zjh4E7Lw090f31T3wPuppA==

`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype="base64", line_length=64, bytes=240)
`pragma protect data_block
nmt5u7gVZVMSGexBbOFMu8On+LK8OKZWypQRXna94i0gmh7FJ4BZ6uSIDYkfXqAR
zS4liTZ8a3VhtNW/MEK7QHif3k6xNmm2UTavM633B2LiX5MhmnyLDY+w0LEsS6cn
Zy4EbDjTseIcktydO+/P4fsAayZzoo0vM3CxqyoccSta8CfFtGIICHYsB7I3+141
ZYcV9/joQlrRA+l+kSkDp5MBk2Q2L+iIu3SIHkkGAk87ooUC7DrKj7kYGpV7MAOS
DiO8VAt3S5zkrUP5t9ibXIYpUH72bIi6CQRxg3fiqE8WM/D6GPjunaOW4F2ZizbQ

`pragma protect end_protected
endmodule



module SB_IO (
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Lattice Semiconductor Corporation"
`pragma protect author_info="Lattice Semiconductor Corporation"
`pragma protect encrypt_agent="Radiant encrypt_hdl"
`pragma protect encrypt_agent_info="Radiant encrypt_hdl Version 1.0"

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP15_1"
`pragma protect key_method="rsa"
`pragma protect key_block
fS6v3qgulmgNE78YnYwI7Sx4E64olqqROJ/Rhb3i1Fq3wXQPtwEbOaCWGi8W+TWt
LxQdbqcFNn6iB6i/jOeoa3yWaahimQDlYPpVi3efPH4iA4vH9uP7/6HNXqBs+yCJ
6A2WfIzt4gmGMrpKYKr2hhZ9ZV3bNkLmcdPAu2nAne8X8+2uJTciMeUYE1d18iab
DcSZm3pg3aX567kVe/zEl+erOsEeD0ElzcKpPVwIXHOtaab0ePrmPo8zmvrJr5+4
0bDh3rIcGK78b363dx7fJ+ThEhgF0rCmaEyeyZdxrF7ITd8K9LTKC0mAiHZ2NUjS
8j78Rwa1w6UyehdIXJi8LA==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
wUXZResLKPx1RKsLH/CaWBLTvwRcNK8JhPBhWN8QuV0RrAmDq6NWaV6CWbyj2fHa
FYj3mQKKUnDIRk4jwQCNIfM/uc5qLCh/RD+p5n+5KZFaCPAdvrRg0N0HiZFyinqV
umGOx87UkpqVznbD0DMsOo6dnSPnEeJmjE3EiaZt4nMftcUumjVZMbV8G1s9ENIn
vamLyEQO9P2GUKlAn7FanKVf/GLxTJOpFYhtEQPZjjxZmsd+0S6jnn3IASUfya9G
39EQfTMJreF24HaL7d6GOcx/LMBBR7GjIwp3FgJqtNHG2gdsnTMvfViZLodKkBMM
4UsjcaMnIHTWa+RRYxrqBg==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-2"
`pragma protect key_method="rsa"
`pragma protect key_block
bQLNwVJBQXawebwYAXbknLLwtJnXVD3pc59NmT/DimI1M3AXQIILfR4VV8dvAwvJ
YP8UcjJhVrNaDHeqwu3y4mmwmIrvZc/5kmGsuNH0mk011sgw9czLZ1r5H6kZ4YKH
M8cCi+/j67xv0XFC3R/KBVQvdtKFmlOzdrJRTVPAKAUY0W6HRXh6kTml6dp35vek
81o7hD4qAqrkZc5vs3SvNx6ccAQ7zcT2N/Lb46ojcGEYrPX730h4aF7OKeWQ47S2
HqXLneGCixP/O2+CYEI+PUon2XJ/jtUg917tvSAgmPz+qr/e6ZQRrAkTds2w3xOz
Bhp99OlVnMbak2jHiJb8Vw==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=128)
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect key_block
g9MBwv4rkxRnLHywvJG7PvpscVyDG6ta3MTisuRxUB2KQ6v0HMqc6Z5eGvNCKxHf
4h4e57GfxWe9lmybPC3Im4w1HysJE5LbdDbZ0CJL+PMoxcxH2sJf4XVyRRdI8km5
d14umNRHiKr+DcAX3b9IBm8WOc4JZ7hLm3rc8NYIlno=

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Aldec"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect key_method="rsa"
`pragma protect key_block
FILD/+U9aJL3jnKb/8pkb8pKvc4AgdCkktjvKYZRSNmhoxCcp2KVPWgVLpvve/6t
JhpMuGw70vq9Iv1GYL01z2iG+5mnfQvyTqMTegchXisFJ7jwH/YbDzAWjeF31QbX
If5BnhwNyi9m01g4KSHolm/IxjejGA4ja+YiLT7i2/eerB5aKYGbxHmMY6BTK4Cl
CGPW7T9m+nMyOKAFtUK24yAJ9XTcPeWFtpxKvNk7iRYi/tBRCyqHAgYDrYXYLiL4
oYEjl7h9k0TRuK9aellpOMAcoh4aLvXAP7TaRP2jQDzu+no6y3Hsowb9kKx25fAC
U8pfPdKwlji56hQ4Bj1m5g==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect key_method="rsa"
`pragma protect key_block
NAB/h4QOn6l8Z1+hScB/1kom3aZ5HIx2ChZJHiaIk0sHMN0pBbR9fXwRMLAo2dMA
uitwZisflW/njBYs0KJ70MFMuionbCh13Mg9Xii34UcnLYMDR1DaPYl0AwJOi326
l2tIE44UeYNuxPeWG9Ed4JUGDU1HgHpRAmSeNTDDEi3RfBrB2Mqd25Mr1UOHvL7g
hnbmuZAIfDcT9QLEtngdEDz7vs/zrp1Kn8kFm+IB9NJ3P7yyHcIckZaC4fKVRplE
lzGhmI8aGrzXxUzaUS95eEKWCDs14qKUKxPb+xHorZtmSnFBezWSC3GpSRDd+NUR
LEqRqGVqosewem491U1zxQ==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Lattice Semiconductor"
`pragma protect key_keyname="LSCC_RADIANT_1"
`pragma protect key_method="rsa"
`pragma protect key_block
oyXzSD7XOV63S3wK49SwlScFyTt0ugqjZQvJkYfaj9YMxr5kukpDt3HxTUnRe0ag
2Au70SHU47SmXRPKUCR8SxEdnEvDzjhl5BSkNCFxZLf8sLf0o6sNPmj5y3kSrkpq
IdU9rIHW2AISpo0wSbzM0yd4ANzbt7byAk6zcAKanLUEYH8rmCYHYsY31YJ3Hhmq
mqJWM++nN5OoVM9gxvyJe9sBhl7um2tmLehNOl/7Q0l/a0c6QbhSxN6RYyPaHw2A
rDTPCbyAYz2lzcoUlQgNokcGdPfxGgB6tr/sUarxYp63Gdniw6TZyACGAqbjAzRr
AWy3hi14oOJw63PMfszdHg==

`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype="base64", line_length=64, bytes=832)
`pragma protect data_block
GqANh7SX2edS8sYDsJBS9ICbkzqnbe2RXmShhdljeQTI3gr4wPCxGyxx15fGUi/C
cQ8NxEiHPNWOJsFUkCGzcaTWqc4UtCdtVDrVd+eRiVyT6YgtCmgKBPwqv4oJ7T0v
YktEa+vtFsMpv/sEwpLxKwVSAJhr+0Q/QjPy5KaJe6BmP8Rwv6LOs8jQ8yMcU06e
KolL+3RcCBpDuUxaaZzBHRLdgmChrKVK4xBGIZq5y+O7XmJm1cvg8v5qeqNFToga
M4eNYpD8edUml1mDxDhBLpbGcCrDN45eZWgsfgLs2khXKU6EYH9tMKV1GvnIotU2
tYU20UMy/09yTf7n3srtCGE9e2Y+DNkQNAvtq0GTnGDhHouKSDmg88pCPGEY8i9r
CnoQTLqcwvl58Z5g8SoGOotLGvklhGi1PsJcry2gLtTs9SqJ1Asy73xQFNWK/duW
wSTsbGe1qdi4D+nXkSt4QSWpI1SyflMOcCfgUamMn6LJpcgEBVuOCPHgU9H8DhVM
pyjVaiVHS4RE4ZzxJSfmkGtUjVOez4mwduhn2F1niCptKv8mxBhVTC+1mKqaWe6Z
GcslfZRLjJgXherGVoRQVuAdOGHem/qGGDeGafVPQkBPaSsl0pcng7jH/PxJRnhw
WNSO75XEvt4ko9xqnrUM9MqvxVR+2YQ1ffsW87L4wWkv/eSM22Wuxxu1T4Z1jNvz
I9PdtT/BGwtrB5YMx7z/aQTjFkLY0jHnhteftx2aOnb+m4I/fPQ7hSZsU1RHlbEj
1ZHP9CfehKkacBg5c5PGZUdXYf+d7ylvNBZJWdcx5B6XC/Q9jTSm7iUDWDZ/81b0
n9xNy5UdjjhIhLBRg7wESq1z4oKkQD9tOvoOP76ucaLR4v1T4d81VHc3Aea5+Q1p
XMDhhbRIX8kDSsRV2ZPqhdiuvMsBEHMGN6cH9kRQ7wPIk0B7UOS/9aZG3/G1v5wa
JgVbspiZAqFh97YZvwypaXDFumM5lWn7+upRdbMh5LRIsd2lGzquv5RPI3QCUk9R
aNw4WICAuh9vdCbqZ1joyUTdUctfqXtS9R/BNgZExWzfTvCrK+yJqr1MjohF5t+c
KM4U0AG5dOmzAuPbe9fzcA==

`pragma protect end_protected
endmodule



module SB_LUT4 (O, I0, I1, I2, I3);
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Lattice Semiconductor Corporation"
`pragma protect author_info="Lattice Semiconductor Corporation"
`pragma protect encrypt_agent="Radiant encrypt_hdl"
`pragma protect encrypt_agent_info="Radiant encrypt_hdl Version 1.0"

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP15_1"
`pragma protect key_method="rsa"
`pragma protect key_block
THoEDJP2GVdnh4Dr4ShhvIMcUHYiR8emJD0AK47/AWdQuH2XQgZnY4ttQBI+ABAW
rfA0glWoy5tSLwFOfzxjrjbY/xwnQT6HfE2rcijDdyI5OTUx+iZORsAalCTtlzuz
2gx5z2971cZW7dv4a2gCUO2mo/k7cmCmNSuks9Fr7XFHQJxuiIxY6bjiTDIR9y9b
jgZBNlwMPUYtJrVh5c+aTpZD1qjp7+Yjl8i947pnziFckIDaBnm7NYa+QfwIajqN
o1Xla+lI/eNPK/HE6LT5/qSco8KmLC+jHXgWxbqr3SEKfKh3fSK4BEkcSyu/iIdM
V8XgN/lRb+mA6YzUk9Qp3A==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
Par/MvTVoIFteJo2ePuk1prfworso84GOBgCt5bX39qIoo6udWkEb6adr75eEfjB
iCMD0aBo/CNILxrMSkcljBZVQma7x2XYInMWpYlhWFJqTp/82iqe6t/SVAc/cR2v
PAvBOH/GQHO9RHLiwW7JtjA+sQnMtPzRukLc37zqNrmVEFUG3w/tEu5pLPAdOPvl
rupeolXEUsw8/GcbGQRZagPm4niDlLmsn8HeAi8Lwz8BKhFNY9I1r9DGH/4n1OSV
WM39xN40A2ufoOIw149XY1TLLEJi9ZEL8Wl4EO8VCyRZAipxcJ1W0si4VTqUL3Wz
IKzIxRuGIKLWC6isMXdhHQ==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-2"
`pragma protect key_method="rsa"
`pragma protect key_block
Y60ro685iPo1JlzTuCBt5abejhZ7X9m1FfoNPcGlqfGIJoP2eGJ2tgFCGYfrHesp
QeSIH+Ts3FFX9B0gBvzEeCzIWdfzqlfvi8MJybhE/uQzqS5EFZexJ2e9WlM8G6a1
ZzJ4g8/n74/Hy42p/JQRChKqc+cCAc4x5ap+JTvM10OkbKK79IQnLORqJsTswzIs
tB1pTDwM2f9gGUZQmeMNo4S1xYzjO0N7I8/udoCLtGQI06TmK4+zeSIcXxOwH0Ph
AVv8p91nbG8KZqyw3tPPPtsGi6vENb24LM/Kd/kzQYsMaFyA60LJLiFAT4Vk+J1h
rlQuSsj8OgwnCmLOWW5mqQ==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=128)
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect key_block
EcO/A6P30p55o8iXHRa+dx8NHt7x6lt8DvFEzLm0anJXoCalRgtk00FN/82pjWbP
P1f7pUetD/kcoCtqE6I1GB72aqcDBqvVyqHMljyK5GF21+k6iVWHRsrYcvvRVIiq
BroHofPrSHVELn8b8a7RrvGlkEXDMt/3hGtFG/2lIhQ=

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Aldec"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect key_method="rsa"
`pragma protect key_block
Eecche5XT95QXb3ejFdBF1gVlIS/JegCiTeF6r4i1wzmEJCDdxKlqXueabbRcf2x
1JzEtMMRQDS0yeTgl1WCb2rI/y8qUJFhBRkr8au9h9kFSb4BJmRpUt/8+McTE6fq
eZXkWlBn58+GPYME6CDPgEMqVELiD/Bgp+GQX8ftdk2AQZFQrPfv9mPTtiuUqUdG
hLgsX8GdagRWsJq7Ueg7M8s+bepvC+nU37TNkGiWHqM7ChnLDUyjlNEtMNG8AjAm
jy2g5F0uN058eGPdq3UKQ7qNBH5LRL872/9ZZqLLHgrgCGI8aiFfBSNVUbwBR+T4
wFQVwAhCHW/rNwAGBP+31g==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect key_method="rsa"
`pragma protect key_block
WrDUNzuu7I3xGwvb8wSGZCsuB8icm9uUspFe8WTLdlmfWZhypZMERY6RC5mzljy3
PYHmkbdlS4amnE3DznxtrNJhfa0GOP3dDuZmr5sBJzeY/Uqkz7Vv2gzdI37tgVBt
yl29BcPixmcpzGRQ8JjRfBNRhJZfMbIjoFy2TPoyIgFk3hyYRKUPAM6dNRRBGBh9
1qyYlbYV1r34932bvUr7pyfPlyhpH5Ugo6SJaJVOcIReDl7CxtkMl+AyUWmq8FJP
OSga9B9Ph1wzvKx3fVa9vJPy1O7k1iIC6NmFeiPBcB92DhTsNrQyAam74MZv2FGc
jELzT42iF7x7fk34gg5xVA==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Lattice Semiconductor"
`pragma protect key_keyname="LSCC_RADIANT_1"
`pragma protect key_method="rsa"
`pragma protect key_block
DUlrZnxvrTT7gtvh3rAwHJZ59mNgk8aRl4omwAwHKNkr1BVzr0/ivvY1ZGce+ip7
CWYq6diprovxWaxkn3umNF5XCPiEl93f1TKl0+8D/jmImdq/y/GX75zphbw6+OjU
ABoyXEVkZ1AAXIQBnMCUMGsZbuI3FnOJ43K3qJMknQFs6Na/LpaK3FR087kS04dm
1AQ8y0t2BDygdPAaKDw645y4A3GRRXcb/cyRDbsKEhOnO398OsgXny9p6uAn2qFV
1dOiAwoxt2quQ0H2Q+qvWOixPPKkNRl8tbkZWWDTUWPNIZ6rHCVP+ZFpYZ+1fBXh
9d4DPvC04UK3BDWnm5cabw==

`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype="base64", line_length=64, bytes=176)
`pragma protect data_block
ZKsHBjE0GaBea+MeQM5nOlA2U2JgI7DDpYNrbGo09lJA4xeFnj0y8ua+yLQZa2sQ
ZchrPFPJcKa77pA7vackcpcFjyPbc3lb8YvC5udmF/LboGkELk8dOZj9nKuNu/Zr
Ndr/AMuF8mhuP0pdw1O6/+uaSUaUPMOdLVoSZyOYSFdM0xb+49pQRK7TrJ93NNfP
505jXM4Vnn4yOkstJ0IJGrARx/rxmLINzQqNBV6X7jA=

`pragma protect end_protected
endmodule



module SB_MAC16 (
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Lattice Semiconductor Corporation"
`pragma protect author_info="Lattice Semiconductor Corporation"
`pragma protect encrypt_agent="Radiant encrypt_hdl"
`pragma protect encrypt_agent_info="Radiant encrypt_hdl Version 1.0"

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP15_1"
`pragma protect key_method="rsa"
`pragma protect key_block
TRNZSnbohaSxhh+ndIQ1e5lIXzpIbkakytc8Tzm4igoTTYkfpPWy6k5aKmc4MhAQ
xgzfLvftS9uqWECnB//UR9fCj6eZkV71eXJImmdIHq5xBtYWwM9lgMxGzLwJ01OQ
JzG5B6s9/azBsQJ5vcX8EsH3DVkxTluIjPk3ccRw93BmMW39VOsm+dq82CZiTlmx
cXKDZ8g0SRQV+C/4WFfEqnkTUeng1FJeSYebaUing19isaFQ6iGI7fmjY7woYr7R
pGMVXQeCSfoUj5lvpBYFHzstdSb/f5BSisjlD1ylDd9gtb1Sq/cCBwT3WwnXUU9a
BqMDA+K4Z0BA7JPGI0prGA==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
e3WdIQFuNpwShUDEtuE5k9fCyBrqKp9YKWWbnUd9iZdYiLH0jV78gS6EtN7JILZ9
t8OTGDkLyEhOwnJ6xw1i4+I4prRqTHMJUKyZlZQv8R/IHSTkBPZXYHFA+xBAR0cf
KlouFGtSVO2SnnPuqu2N4DbugJ6bxbO8csZWyWYVOQ11bRXFcXZanimEIPZUwdPB
xP0AvnRypss/G1buRIdDgHf+7TeJ8XPQ7PUgHycwCJrpuRz5ZXrzuIGtuHkUyUOo
4bAnVDt39L4g6NIRhA8cksJ7KFPzVgMWmiQLElBEz0CUe7HZaFPIjylgpJeRXqal
YyOiTVtC/fu/WG6dCYgw3A==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-2"
`pragma protect key_method="rsa"
`pragma protect key_block
RqcEdOFS7OsQwahzIkXYLAKcnthUAblmRjSc+AFTb48/mLHUedekh3CXUtja1k+l
+UvnFic0j4PF19K0LACPp3SvDXv9VBq4V5WcDuYw2hwb3bss3y1HAl+D/5LzNMF9
IPdZDmXADTBApmIpx4fzadabJFef/T4xcAtZmOuYUiQHZONvII9c34v6wpY6YDkI
mPtscqhGez11Jri4WB7Y6Bz2M/hXKkmtQYMrHTl17B0WMZii+v8telIv1NPF9wh8
vNRiXAd7ECMXEQmiOspGC9KmMfcA8PTVWKhfHNwUj64Xb7eUmA57Hl9V5BwY4vf6
64L9yvurpgAgwh0TcZr8Dw==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=128)
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect key_block
BRVqOv9llkv+6B12h+2z8M9jDpzD+d9Kl93QwpAWZTnsIILKJjGetyKUDe4FXCoA
Mbek98blK/qWr0almZbl8U+Rd0AmOW0xNXXb2/musxslcflW3gZG8mKUcvUhDR77
uXwms7q4awo+10DF2IppZVINmTKIFgo5+ApIKyLP6f8=

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Aldec"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect key_method="rsa"
`pragma protect key_block
AcDsojSgz/m/yjsZQbGYPkQynSxte3TD31owd5iwKAFpDwsjekHr0y+jSuTmv6u2
GgCKPppeEbFTEEXv45KgFRPqMbleOuc5KU5A562UnDxF2Lm6Cq/S/L3WiSASKSDx
1nIXprpDoLKA7/KXdZMqACREQy7bSkoPUXYwVCay0vY9g75wqtdYS2I5noMuJk8f
SZ2UEAzyskxl2l8h/CXXpGJw6pwZSACtTRvyG3aHepMopFsEQ+EnqCdnGcFaRguk
zUBFQ+YaK4JKElzY2msM8dKLYnSb0s4UHeKG9ZVSy+O7dcAvOUwm1KFGHYdHciHG
ACraVX7Ip5DDL/nniKMJLg==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect key_method="rsa"
`pragma protect key_block
S+v6ZBCZWNUFXM3+psKWpHhK4toU2wYmpzxMkhS3GFy3C/xARpsWbXeufeFALkgF
C48Ggu4oWvOJaCMiI2s+1Adh5OQtr+su+hzbzOyAnQDxfrw7PNK7ge3ywSnpENn1
gws2EhFTIBls+RILSBpBaaBsNNrPCCMY3Q71YkMpas8mCZ7w753joWX8suLlYI08
oWc5qnGCb0udyOeG9Q2OZ9NWPtV6V/l4UnCwQ5wCQwBtKsB+Z0B3DHRYGg1MJ5/H
sfiRsSVC65LIgm8Weu+2Wa2VV6nVWICNEjbKnndByxzQfetn6DB1G+dxEehE/reR
CINRz49y/1NtwFw/8TMzgA==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Lattice Semiconductor"
`pragma protect key_keyname="LSCC_RADIANT_1"
`pragma protect key_method="rsa"
`pragma protect key_block
yzGsKipChhIbPNWKso+d1ztWV1HLI7lEsXeY4+E8qfdA99WXVAej2by6n/KA2pn3
oyxm8MFM8Cie21ptAFFzTeIGXt+fsvQ69QXDkB+YZvvlqjv2y0/ufxXb4tiuiG4j
SuQZ6ngh40kJxhdRUbqtWW2I6BqWYoHor2e238D8wjN2OEj+RgJvySkRTSzYNtie
ya0ewDej2PkzK/EKzH1yuJl/HWup/nujM+SXotrGidlNrEcgzX+k6g5eDJ1HR6Zu
wIf9n7U4h0xZru5NNWGpYQwpgOCMb+WfCbiGxNhAW8FfzawW+tkJltHn6oYNHJAe
MYi9QNyxBhUp2Z5HwRIcZg==

`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype="base64", line_length=64, bytes=6992)
`pragma protect data_block
wDquHUw9J9GakR+P0V2Y/dIf+Fq2D2kplIp6X1sljWv0TA/OCRbUlGGMoZxbHl2e
2wIo70lMPPd7Ypu0xK1m7l24/AQy7zD77qQX0699tb4w5jXLioBsSMs1RK2unUL6
6nJYowGteyHwfVaiKS857Ghjh/4twlm5WJGBD5bKGZF6kGztX4ZX/Efrp+X3WalL
aKfBwNffZJAAfXtcpNfupf7xECXYLUdJgpzQTAKzu4OwqGV4FgtuVR74hMgWQUzJ
jrKO8a2is3SWVRKw/fmTKO6yRaC+CfICaGgpPtP295XLyA6Qaz9vniAObJP6oy1A
RSW/Kull0e4SQVkP70jgDPYM66ZLN6n9kl7hHM0fODsCa14V4CxWjh9rDo+zXSJl
voaaeSc0DOvVbNXk7BuLhbmoWyIcJBhiQkZSrn7NipvWDJi3/2O7rHHD7kj+BZrX
OlA595/2caWM+E4yYfXVsZHhiHOBvBHo3e2OB0p2xQejESQL86sFneYqSw7qph0q
MEM/oK5XIDoOofzajk0Pejdc/htaczTZEWnEz0VxXurSRXSYQdwkfuekkwkB1Mv0
aKxHSyawfDSEymw9ZO9qKca2H7TWU8QvRmtN8NqQa3KrvE+aAs6aRQj3qlyWkp+J
tI+P3waK9IqNkZKjwGuL/Doyii0U79IPCrRP5oxS8oMcr3KW/N44ua9i9q6DX30A
S6w7SIEHEtzWnbVgqpqfjPBuSeQGWmtHIn1vSFph4FFOyMtVz3U80Y1thHhvAhTg
YqSmpfWSomG3ayvSRUrf6q0Eh1XfcnXy8IeFVPug+b2YqD8k9e1hqBPpyg6f3lUt
D+cKuNap0xzu5eG5UW9hITCbBCxJ45AGS3Ey67P6g5Hs+/w5eiExeLoH9tHmUviK
/0nY0qIMRixV0pUTrFlXBBC3MhoWTvJimBv6VdiL/t5AxQmxab8oJNqAzfwJQYVK
Es2ie7b6GpXXYcpmhbHCaFlyFUS7YVEofNLlYv36QYKDBoi1JXYyvaFuTUySkEJm
NCWbH/xiQSIveFiQZVmRvPo1UEqA2veiI+ezKxdf9OditU5HqyGIKQV+pI2yB9b0
5qOrAs4YPohKCPoDNTaph+lWmOQXYwn6tF/dxfZ9jBErAxSN1nR99+99N/UNCf/R
ef5qv3Ra2pmVoXbvwNn7lavC8i6RA6mUVgpjLeubaVD/ZmuiQfhBBQjqTD2P1Agg
Uj/vf1ZSjt00+DJJsRrJfSvfSQbT3WrMj5gI2q/UeOEYC8CKCcIIiUPMm/ifbrp1
YW5o766xSUvx0L5Sk85AtExyNqeb1Vrw+T5ZZhQSazS3tqndHrC677n/hM17cUt4
oD7w+TlDQGS3IGiA21DCtCQxAorRSxy3Txmez5Y/wjQflKtKgArTzk861RvWYj1D
pawBgBkTGzt8Kfy5/Hs+q2cKs7fxU+fbdEERZ4VM+ch1aRDEg8rf15xCZwWcQ50q
rgWEqJi9NnuyKmdHVIRQok4+XcGukKLRJv53ivUwm7RPF72TEX7RNFvyrYMKbEl1
M0X9QOXhIZ/2bzgfwxHcw1blGuCiVq3Y9W7ckkihaaYHORxUcnYh2i8PK2NS0cZg
tcS1AQbn53QUKSho8x2RLCLeVFTuOD4MzJFVpRTP9lsqA1yKZMKqvPfgyseA42Cj
aWweZNll8k59lyArxJjQBiUmQiy5XdmM20TnkmVU5f2vmzWGK5uxKmIqysNvcmKS
511GDYYvyyIkMqcX7G8y/TqF2Hyy54K5qKnulghdzFzZOvsGP42pOhJjoDeGbStA
sEy0E/R4BCr3BgDFBn0UGnsBswpjF/guJZE35PeReRyoNenaR7KLEY+BavYjpWnu
GHZSPs8JLjTrY0Zc8iu9vL3OVhC83Dn9qPsdCKUVd6b/kVbNkd74c3AEZzwelLss
Sb6pHOZYS5fdCmyPC2/Qq7hEBC1+12zbSx+9iKyQ7Uw1KovqFulTdnp+kB2b8hdX
p1qnZ74heuL+QXs3WzPeAnzss6P0BGqnPbkewgmUXSG3iRgLgVl/KhFIDePpYU7B
1scfTa9Lr/72WlRmWIcxI0wdn4N9S5kDjTfOS34XIwGkcpDGwzPI1lKriYiLvTt1
00/Kyp72KHaIMgcjsIAsl6Qk5vjFDepAt9m9Mp5DHOCIhkyAGQFhf7CwhNHahurE
ZDnIHGZjUR2spZOFEgVYo7Lgr4t7N9aL83HvZRB3NFB33XazmnPmGSvbIrCWrtMw
1gIMDjorL64LlcXYdGHMOdO7Itsz58opHq/r5AJ1s3/13ndMFOZEMLkIUzRZyYV7
gomBWc48NEC2XVIzWzcDHxaxGansL6G9S1Edwla9wRO6bDQ8a+P78KH8FBLav/7M
XUgbtIhiUOZ8gNs31IGKJ7QTiZ/TkbD5n8J2yhfpzsR24xL/psxk15v3vEqG25vr
+rL4jKHBT0zK9Dm7LpRRClAFAg9AVMB12jrO7m4zsd00io37j7R+0oviLUt+ywcY
dEYhQ6EEr7qOuAvbQB7QcO8Sb55qDbmini+AhdSBrCKUoJ8pQhUtIsTdaGrnxg3d
KKuGGmKLhgjIOF6cKzhsk5aPF1Zg22n0S0rTnUKnZqj1ar5ZO8oYs4p5sUvM+n8u
sPgzcvdRSa0C2dvqE5A3p22bdHDOFdA++7rv33k7ByIOLJC3a2qye3DrxkOUKbfH
RcuNgrEFqH+4JlHMNRzIE35vsY+nOv8yEDFthDMIap1SaZNjLRvkZqcA2u/LHY+F
k47ua7AuaymqkP548k0kEmqG2vNg7Zec76rdGKmNeJt/qcjas64QmHTIMtqbotqN
vBCqUf1czgX5sgWu58jjLGY8IhGzwUH/6UmGUUyTVdoTIKmiDwqUZFztwqMI/2ar
zW4f6CWy0mxUIaM3+iKOA/36NlcruD3XBCAgMIKWhnvPtpAwgLjv+ZEzkuO1QaWY
vtKq1dd3CM70kstB3jQQBVqnZoY4ZNI68o4Cj/3cXOtEYN32C+kdwHyO7WyG1u2M
4hNxv3WrWd4sr8pf62BZUuamqTVzR6y7QOnWS8qqR4mBHGXcJFpWZaBhq3vU21WW
hAI9S2aqkvx2JKhQoQ2WaGilZDjR2LkDs8xuaVGaRWcjAS8DwuJl4IQ++VMYyu9x
2VWTOBUiVBOMmO8BX5Jn4rDGaGDLzCDPIS+0b1v7vNNonbBYldrw7O/ZSVUXsYdO
xsidFQaoMEw/DnNta+FWpcvSHMTIgWaCzRK6R6l2B/yKzWdabO3atF/XJAEwje5Y
qE6e0K6lDl+8q8Mltf8TxAG2q5NXbFLyd3Fd97MIUQ0aS/iOm5ZPlO2daVNkC7RQ
DVMJ2PdBy9D63ZQssjRRfWjg9dRjkusM3DZJoDvtmfrOap+12zWHUrIuNh3uTUDF
f24FNPRb7FFxRZq8WUJCUSZOIiCp2GF7iX/Ff2pGc15kNLlqay7kkJVGAu721x6m
UXiaGpkqhM+bqOHpbisQ3znlIAmMFql+eOdUZ5ats4gXVLLdFyKjX+5ut4U3AyHu
TFqqGjzs5LjOGzkDG9nBQP6yYq+oiz6WR1DOzIgOVImQWDVliQeV6OXXlCjAzUWs
zxxYqdZUL2gXXuA5UqS13NZoT/BBcoM8lSDOOZM1RrWC9CdE38a/j40kvTrLOknd
CAz1mJypIFHOjnx8f2dTm71TNNWJw1ErRbf9dJ0Mp9vSPEiAWHntpP9UHgYMSpXa
HT7nkU/G26RKPMJf6XObsFBhfEej5HFYwBuliFsCr0NVkq9n5adpR1H4+CMI3LV0
E870dqv5/tgkfAOCt3kA8+g0201esSvNQcqUPgzU87d7toowm8yZVqpuEdhf72UA
ZVNcEQ8xlAuGkZqYNjq9Hr7WO04LcC1SIlt8fhJm7/0RoeYo2eBdLcPMbiDI/lN1
HRV56FrtTteLlPrXCyiTmr6VAKRheljmmcsSkDIUB/RNBGsasak7U4xo4xdPEPHg
Qbq7ARmYMSLLxU7FAO/kmHytduoXuMhQDyJrvP86DxMKqWVGqxUy4RDQVgiRCfoI
IS7dOBX9UJBUmCE76/AXvwom302rP7BPHA26C4Vdh0Rbps/XVkOQ5Bsyn0m8GVAk
ohBpBo3PwMeinpTXGZ4IVi4m7wp3GnTiF8YxKfP4hT3kEc+wyY1VlNnbIikKxmZw
F8AZFJ3mX9uCf82A1VOJ1aRwBuQ3rP2I0BdoomBEt0Y/Ovq7NEomwBX8y71AfLyC
vyHfp+v5xQ08oCHlPb1NNC0mu0+t3q9rPIA3530L3S4bLReDoEE1PAsn555fK3nR
d2pf6CsAVBVXB75QBEVu08V7FabEOUoSPs6aft/BXRC2BDYqt2tqchnd0rOnZwXW
pldWulsIAtEi5RrNsu/c2pBH+IbXjfRcml1IVNFeKIFuqhAyqWVqfqiDxCJ6K8JA
jowbNK+dczmqLxNnBPjbeleApIwtNumdoi76bmF/rLHWIRcTwtlRbpybAnQ39cv9
Mok1YQPrji6PrZSDiylXIBQn86JxarM4nJyg/z2bESlZbvKjzxtwra64xelcwmkv
MLRDDNUIQeIk7zugihcTCrRMBI61vqOejA4FlhR3RvqdcptdJvARW+Gz1YoT7GnR
NMrkdOLj/VunhwUdbyDO2Nf6lP2TuenRThA/7Rkfe1qGeJHR8r7YOcnxyUhfRI9Y
E9n9r4hRSA1mgAOjD1q5PSDzEhsyUtDWor7Jvz5W+kFiGwfbQDNJHYicWqD0R+Qu
FHhScZqXtvA/S3L7SkxX9qkLBneyPLtv1JRWTq71+0uOUN4xdIN5Y73tGVOaYXuD
cAWfdxbhKQI8nYS86pY6Byk+q2dXVUcQml0QIJfKFcl02vryi1gFnRInNAhM/5rf
ZWJQKaqdRoDAj4e4Ha3zruWHdVw15PO+tKu/fVseW67TgAPgKSsBtenKHipPs5vH
OJh9GCI2r0GxYaT1ne3QSUSv2BventLULI6wa2wWXRe6K1BZOoQmWFz6XkEpfAmB
ArUA4TNvETgspxwjDY0zlYmWK2t8dTs5T5C8GVBAEamCa3DOPx8lUbIDpgioHIh2
WnIqBFk8nIGnLQOI7ZPa08j/QGS874GrhFXe5Mo3WTiBQ/ybxNE7ac3F3BCpX6jh
RwgU3tM7NGecRwdZ7LUGWkJWl60WXpMqm8v+qBs6vb2E0m1m940bVFK2Ch5V7qWM
C575P53KOsVJsYz3REQzSCKHCtMvnDg/lY+Vr4y8ZXdxylt3r+yLIk9i2W1KJu8U
i5iS0xnLaI6+IL92zEEMUBB57dxqI52fS9FeeFxmGR9dbszNKeAUfplu4jJK3YqJ
ryFeXVHzLQOzc0pdqV5kEbxvOn0auM9YtDz3lbD2BQKYLuah+lWzyPHPp/fyxyrz
gdw3hzM5039iDTWLVoOpwBc8zWASYkxjkhR+dG+ZyBkHYJT1tzsP/Pa95Geq7nbR
7PahCInuMLsmApVChNMk7t6/pbfTmsP/GAyqVZhRLB7v9KtbubVzjwtVdM+24rUA
cv64mxkAIOJ+YS1ffm8YxI2P1FZ3igM4MN0voD1UEMuCTJK1mQDMuIenn2xsFu3D
MhK5TOF+1TyZNQIUvNjVgPqXPlL1pJhag/9iQ1MEUcxGftx2FC5jqkvCP+EMWFy/
TsM0VWzVHRuFltx0kRUHeHoF1v3oAyx0wJC8H1pyZXoMokxvjFvDnA6ZweOg+oVe
pQMUfWuKilgfwajo+m568XYRAZRcQAf2IozYbsxg+1+/ZiPLHiewo5vTLvVrX4Cw
vCLN5EKz4Ns1b70E/G/Q+634xAY31fKHddCoA03Tdf6/FXcIm/+XABREzpgDoiN6
+nxKAnn3q7jAbjjTmmnXakzHFbUvTa0uBFK0gcwUdJ0tVPoqZLrJwwuXIpPj18fQ
arGhSCWW67e1gTah6XqQ4YFT3HAMis5ki3Hm+hMO2gb7bxxTEmhJWPWu74jS/LCF
8nFFN+Nwgafev3GcTpFISRRd0NZvXU3H/mW5lk+LngxGEr9CcX52lFj5Hd5bIZqW
ne1iHmCWfx02eGQmT2G8qH7DzBH0H/K0DdUKyeNXLqgCaWrRObAt1zAK7HfCzOl7
wbAZkaxSmD+Tl2ArU31KV64u1s9034QjMHJ632sFoqOPbXOmEgSeIpjyhnjpi3ZG
7pEEdq+ndYvrNL9rskHDBII4Va8of+kN4x1RUxkKmleJocPM4i+GCTuY98eerZfD
N1UC9c9fJsexq8JxEDsIT6X62Yy3efh71bp374kLi/1KVDxjiQxKgCT0H945AD/y
krsx1l1aqihLm6rsoXjz05qNI24EMg9CLf4EK5136rg4Klqmks0YNrDXQ+63CNZ4
QclXhkt9+ryUf4gNYI0LZO+FWbqwsU21fzAjr+IZLsdxyqEP4k3u4NiKvFQJb4TV
Nfy7eEv7hKNBd8I6LGuo2HhE/AAjz/xsXDCL8qrstpmCWMO4OyKebf0pykQJshc2
JSz5rg1z5SMcH66hUulaBDi44NlT4ha4tHIMwVWKpDRVBa4IydDEml0ktS7OSlSO
/PgzfiAFPCJGXH7mHGjqQoaLHspesQ1loI3LQREAk1oWAhAO05XuD2IbWcYVL1yK
xElvoF6c4EV+RiIIz4B1/jyHpLaMtg+sOdGcIFW4m4DrbD0HjmyobRd3cGLIJky8
JahUuRT6wZ4mdgHLvtmjpA6feiufUbi7sU4dfQf7yAK9quJgWjB7WcMtz91iHb/K
r5gbWo3IBMEp5dEY9d72kMk638FAwB/Wed08j8aT3sWbeCpCpd0ETWpggH+OqZYm
4yT94BtK3kDregWUfE1JnCnEL+j1++39KKdBfG195YidYfp9lLYhLTREdKgynIBA
T/baSGd27z1urbmh5RdCxAgI4oafeTRGBr92+KW0KxQXA70m65t5xqXyo425Rmyt
8NUkR+z6GFGVAFWDiuUy8XPtWYMMXapXyTr4RVrHmcmlG8aNK+82fUzdMhIDtSDY
FynvRdrCS+xtspnPpTF92PF2B3E5V52Ehe4ZDJjXWR9gOZZ89+ISczMzoLwnNVJB
P3Z+fqouJDWU7yKllkb9vAAhS34drr9gGEBvUXnbvZmMBX9hlnw8LbMO2VURCXql
tevemSQOIOdwuk6gWJ8eR21vOa9joUUq0LYX2WtF/1h5nL39/plXEY7OcM31oVMN
7uHM4fjM/GajNJGt4bKlnGhNobVhE8MDx05+JTU9ByOMihB4duLmTmq+5eOxlo5j
koU4T4rOE/Yh8euubezGO9NcJjHfBTYNk9/W3o7/bdBRYhs18hZ47MsxJNOtypUt
aG2hW5oZMRtE6+bm01E0bNTXtkdaEvj639suKqoqwtGa5KYvMxoK84/32dtsRmo2
bkH5O00taQSALuX6eMS+mPzYq9KcX03LucNHYfl9GA3PFuB53kRVmXi86dHodfes
Be1w4umsgEsZ6MXGrkgYR+eR15AaurXGoPwbU5D2fpsU3zndOxgXWoY4R4SLAfTA
TstLpywJw6PUU3m0GhMl/MjNEy23kAxnv5/6zL/IxcLrOX45r8ALDe5L7/gDf64W
YeAz0ZVALfdBfWJzQnMeDg6bkNFMXPrWcu/M4A7r4F7XwoDU2X9cALrWjAs/rWla
sYkNrAKXVKlvhqJGice2vsTelZVpp/ylC/V7VbpQ2BUSUYkIWtvj7JJLPZqHUEoK
hk2jlY4AHRQc9jt4Iw+dDQKCVIZoLHjRE2h0s1D7pUnGxqiUuQW3bXOlEEn6ePr1
TQNu6H0T+iEArIHfqsjYGkmx4vM+6/Chop+BsH8XjMDuG9qZhCv1vx3bJwFEZHG6
qpYre6kZnBEnq55hzaBEBBW9h/dlzhrlCZUCZYBupXOyXSKDLbDS1dGEOvxTJECd
tfGdpvdwtteQxlHYau+XOZkPP4JXIIrXx3oW0FUYs8P9BhW6IUJw6waa1S/4TOBa
ffzvjLlInX5+umFmThd69TjKrIv+jiTyWg6FtqkVwEFbmSySOCXzFrwu8OYjllbm
FZEsia/SY8e7IDSzELtOpr5ds4OGMWFMnCJflvs2DWdzRTncj3a8SeiE2iW7Cl6v
5ECuitkZ/p6e4msJM6oL3XlgKF2kA7sKSAum6cWCmMY0XePfIvvXsVxbfhUsZFUv
p0fOfbPldw+4DuwpWrZX5lBgvCEuIvcTxO+vGpiGmBxJl8xrAe24O+E/HSbm6t+A
WL6YnHN0NngberLJhlU+TunaH4QIECTx7LG6F6jt6XtLfBcbQ8cPy/vZLKyXquck
TFSeXdpz6PC9FSj/cqJIhuTYUHvNi5n/kRjnllQlW+xw6oy6Ze6bf8yd2Fm9MLSb
5xtclJTstxkwAC+B6rh+IomDdjnPB7sGYfU6Nqvoxol9dep4sPppGrPpJ8CZrhh+
sjUh46nEtcHhJvstG89WpF6MoBsQd2Flq+EWTml5dLTO0kAVwUUiX5RY/mFxI2hp
cAuPp61UiZ8mG07vNceU89x5uhbRmobgtSWf16nMSFSmcV98fKBVCi1ghcOboZAa
oWxrwAbD/UuYy5dRNwgT9+M5MlUe1jhywkI4F2ns9ZsCMGtQU9xGiYuvMf8Qly+T
vhreQ4kNQZCoUZ8b+hc/PA7G3JrvDlIoYialnCSM9OUD8Tn7Ryyiq6kfir1yGWsV
PhtKMWdTzrRN+KOqF8cpYgV1ALPTN1ZZYsMEJhOe0XhAar/rhmNU1nERL1orRbKu
5e0GsHFa5HaQzvzfTgmPzKRMmI/L+aJOiI5WU+zQwiXuWTxx8sYD7LdLvDlRXgdq
AIl3XpP4o3IGlcFlV1EIsd7aC8Pdv28HGkHOXymbu9PaiOaAO77s+F8WLfwkszNg
SXmO0eFvr7DoMitopjrC4hO4NaId86ihunQC2QhTAZiqrgSYWHm+XOhDA1YbJNYw
i7ErJT3l0Ei9rm3BLkj7E9+eNkRCjM/sq8Sa9aMRCbvSDQftvGtU64eu8sDB/oZZ
r04Dm+S7vdK7mLwK9r/NZQJ3NAH3hbhZ3FdWfdwF93TOIBFDPHvLfEKxZSEY8OFQ
ShqfqxTubN9mx+PNoEjXqAoUV5hlGqa0+Qlfj2OocZELIqa1c4vjpfmHhrHBKwuw
SW048jNY7tJBKnzESDjGYh9H4PvBefXSHp1AhNNLXMgpzego4fmXzIzOb5NtMcZ+
mkfUE8bGal5GzCcV2WM4wcx6451HqUZ/OXnzheHL0MbH57iMsV71940rcoh8JGCf
iW4PSPNMVkBKL3caoqwcfbtJVrBXGLe/A5Cv3SRyIF20YzaoMfqo6pOAsZg6cm+E
PORukxOJ78sVfaVxcyotH6RlmZ7IzbQwRPAv4p3z8no=

`pragma protect end_protected
endmodule



module SB_RAM1024x4NRNW (RDATA, RCLKN, RCLKE, RE, RADDR, WCLKN, WCLKE, WE, WADDR, WDATA);
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Lattice Semiconductor Corporation"
`pragma protect author_info="Lattice Semiconductor Corporation"
`pragma protect encrypt_agent="Radiant encrypt_hdl"
`pragma protect encrypt_agent_info="Radiant encrypt_hdl Version 1.0"

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP15_1"
`pragma protect key_method="rsa"
`pragma protect key_block
FZ1sfyrzxJTAlAlbDHFqSNaswu4hcicFQamSjRHJbxc+55MZI4bVoWXHyyAEq39q
Uw6djQZvJ8St4l77+DyAjBBIdwYSGBt8u4XuEcp+ciIVWC7JAnNpBipjLbQqnDDN
dw09bpYz6WeC8Ven59xAJ8clc0PzCUCNStsbCJL5l1udoPToN05vnb1ztXFCzQxj
3U0cggRgI7oUENxX4HP2nmBpQ02QNPnPQ+3uGx1wRlzzVNNEeBljHappw+x9Lpk2
fubyENeoDuyYTtZXiaaW9plFSZKQrkru0zHdzFgtP9s11t+uXC2n++x/cHqqemPz
tHGg8BE8YAwo8rn5H72nqQ==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
IL5dkdlTr4LAkfqo7KKzqOrGXaXg0gWzGYyLY8kxkGYKZ2GnrkjiqY3l9XRNcFct
yjd5BupOrN9a6A1MAbW85KgHzdV2aBzzcNZgU/dd7aZ5naTPbV+8Ddd23+QG4CNm
DZmTlYHYGJvaquZSoe3CO2EKIazCATroNJ9qCTK+Ks8t/5qIQPnG5SwaHiK+Zs9f
AUpDBowNBYER9Y1ARR0pQqedxEPJDPxW4ux5M0CJOGm7OPvKCiU60lIYC4ds2qzE
xy3HUkLtXBgnC4GW0huk8pWja2PG7lTYbOhcGuAYQE0ABzDjkRRhEaboPSkAreRm
4AV5Y1Cy8hMVgHRpkMeAjQ==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-2"
`pragma protect key_method="rsa"
`pragma protect key_block
cJcZHZ7K3BMoWnM+j9QySmSTcejq7tu5zGrPCBbNBXMmvSIqaAIjp4f+MJjmEjMM
waoCtnnoApNWlSSyvbKXmGmgEIr284HczTz1hXTHOdwViIH/7PQNSuaP9l0iY5dQ
xyOrHCe5Dgl9ElC+frjpNVg+YrodgnYBUVS7qzBkHE40GXOpKk/axAWd7ZAeTiYu
Rb7KLhGPmpXcXgjrXKUPHAnPXdWkL+mNa5D82HlOV0HechIkgiQJx2oCW9EyTg9/
6LW8QOLGBu1Em4W12Hbr5FN5FveMh9r6KjKm0MxdY8kachEH2IDVdfwEqpMg2Kr+
b4anMtk5s5dNmBorq6v2iw==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=128)
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect key_block
D2X1g+pNZKS6v/yywm/PjUeHoN8Sliq4hZGMkm8hHAj3Zkp1GmZaX8n+4/7o4aEJ
T2bkUvvroWBkjWQafVH4GHZShQBZNh+7E8RoMDpp+wCvrNJyU0QQTbUpibLS3dZS
LDsTyBAS6Yc684vPcB71sP7VeH5akIuGRPuhHJ07Y9o=

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Aldec"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect key_method="rsa"
`pragma protect key_block
ca8v3BmApqay4ldzuT9834ELusjkt1YSUmqQDNOmDTF8OcGnKnhikbjzAhZccKtr
YtzDAxFdu/b9DFeSKDoS7r0gkO6Z2roRYZ6a2JNp4kGZffMs1Ph1G1xKUH3JZOJD
au3SiQ7YoMwRQC9i3ftwlTK/t25tdRxtTW7MQZKKuCft+qrZeR7Lzuymjwn/fgrr
JOcVukn565jImbJkztt7ms/3GFF+6anWhVQjdxVemfQFXEz00ch0xCsvoaGGzPpQ
IKB4VaejLBnnYEzE9+zzXmkcwiTWOu7ehiDnKC8ATwIZbbTEwA1CSvLbyTUhUtqR
wrP26cdnu8h/l8h/us+WEg==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect key_method="rsa"
`pragma protect key_block
KnSvMh9u3yDC0v6DFOMaHXqMI/3tk1yN409bLojYyzTwY3+x58I7FMW1PtMcGTav
+rVqtFHOHJkyfJLNU8h0yqvfXO82uSjQDEzq39plaL1MfTRuH4g8FodxJszGfYP0
6A4dX3Oaek0RV9CUayjv+4PELK1owijrZ5W5KuIYhyna6s6vIsnGTAj/tgi5RUYt
givCbnmeEHi+y6zqVH62v3SjFXbVFUThaiigPhPy4FvvqUhYvhJqKKqfCDQUa3Ix
p9bjupeoep7X0QwpevyDUtO34cGrIeLXd8YQxXbrjzEbbQdkEGSo4gmiTP11Kxpg
MQ5NJXLkw3+BNgEePqEsBg==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Lattice Semiconductor"
`pragma protect key_keyname="LSCC_RADIANT_1"
`pragma protect key_method="rsa"
`pragma protect key_block
WnKwcgLCt/fzVzPvFlZtS6dS0stXhvtTrduCAmaYpuDa2u+yQG1vuzgshBahuDxM
MMyiTfff+CRLHnH+nySf8ByzhxgJ4n5tph3yvo/ez3/KyJ5qID0hqkpm8zfhNwo4
TrQkDvEDKiIWciiykxnLDDiogpKf/Y6nH2lJxmuBf/GUVyLVlZUlCyfOb04tKX37
l7QptVlV++ZQjc9I7uL9Xn2mG53XRpznSU8Ro6HTmTLHb9+kG0oMMw52G/fIY8Kk
3D+yhetH80zk2UiIaItnmD22Y5NblIQrMs+PB9hNrNeN5V71xvahBmhwz0SFWsr3
AYk8LdOducY5GXhO9rcQNg==

`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype="base64", line_length=64, bytes=3952)
`pragma protect data_block
6rX1cB1ZWJ/VUdX1gaoQieb41INa0APYZCpeBBfoh2iZt0QLAq3CqadJRotg7PH5
l1qDfVJ7Qex6HZOAxTQhRn0Nu0rSm7NAD+lFY9hFO+dXqiuiUmvXBqWCP3qYLjO/
GtfUwmmFQvf65UYjDheGDyjAjoP7I6WS9/9jItaAOweAbibVy4VtbaeXyS0dsLyX
BWFWgvozFGCuYMk7ut12y887CJz1ApPKgTtwluVcyIcN1IDts69SsyW7k2jbr2Os
lfgns2XuQuqQH5hNmmlG50HFe5phyhmEZ8umYPOsobqIFu0WgKTy6EdH6LbLlW0e
9dDIj8qcfi4OayMUgGHXCwkKCAk+rXCsPaVIKlirTEgfd0wSgWeLsjKMA8vIMN2Z
eOvShzb7+kzbGHs9vIDIIqgqTqco0y6kI3ZctGSuk4l6jIALhvbXmidMFqAmSmc1
8uqFoxz0hCwmTxwwgpYYXKS5uyhWH0Oz7/WXdg1A1Ls4FNu/Aj0plFmSye9iHnPj
cwQLTOdofD6+nNVh3B0JsyFPq4Fr4RxKZ1AM2vMaKx8Vp93qGdGlezYAGUDaRhL1
wyIMg5eHSoF0t4kCHdEVdVDJEYCAxocx89EeeLGuBXZfUQBwGZWfluzmBY+proHs
Z8RYMmD32Iw38fffCju48KJ87lDZSZ600kLJhFhqRLzTeqLPmtOkx6X5Tn+q0PxG
f1nuKpXYNr8kC/aK/a1rePmsAv5MYRrRiLc5JzLD2g6a5yKevM8EkxRW8j2iIAJp
q3q7PQvdXa9hLyC9TJssvZw/NVuaDlJ4N9Di2vKXqFWR9NhAFk2j9s834A9VJCmC
XubwUzoPH8WExpMeJbeat9aMzw3aaU4t4+I9GYDsu+J8e14qqTjGaZa5uD5e13LA
KSdsFb3A9bYRTO1k+GKPP52rpgj9lIa0ir7rWG10INFI7KBpsXSjCZOSEgpDJwLZ
YZcXif2oSu7r1c+yewsdp/Pzr0bkDAsTB9LoulDnkGOojdqPdMJOJl7pLsX+JLrw
eSuFaltfzwMripzV7JWm2envANkZsetZsHPvWK7OdcIiTsu+FjzxnNZoADQgjuwg
cy0qmXQR5mTf6im6F90KNQ9Ulp9ZfrQnrGAfPi6GiTOFKNPXIym/xV/JltzXnWKv
a3SJQJBSjAmA2I6fA4QAOKD2ZOjsqj/U90qdVwvZQ4C3VPq5sJ9OysTU9Hqxvc1H
fVmSYSHiZ0HlesX/CkwwRFVDWA/rvv0n8OLzhU/hW0Yv7tNJrkf5t23ozSZ5zTy2
dhEZdo3Zx0ZdfbEtVxQ6a539yZXY0prgDQrLI2ltkbUgTvQ05mKuiRuQREM2MZ/v
CmfuTm/+G++koExAcOypJvnO5Cy3LugcjchcFOY92DuKq4+jnSQ6uolSF6kWxk4l
oZWzx9YuMGCx0TIcq+/Jo7wpk1FXqUV+ftXWv3T0WdDQ2LIlMeNnnUgIE12F3ugS
e4+kwM46Wa7drfC/Xwx6vSIxko/icfx0VS0Y61cAZsvT/Z8c43YBxk7X2fdLUdnB
zqEdp38aM8Ok8Qx5+Xlp+IECeMuYoYu3Bt4aLCowikc3S/lueUoGdiK2iDPHpJxd
GSOluBiUl+vErH8XYVxc//HVUN6fLDLNI/crwY6MVjNtsVyD+Ek8ErP+y1KXYMTr
6ssLx9nikZAkay3fwb82dbwxBRZ5cphj0qOuva9SduaAggwnrTsNy3b3eSFRHi86
06FuB5sRsvFmrWA6zNE8Ni8/S+ZZciXag7ySyXppmxwq5W8Z0kuQQo2t6WN40+c1
cCMKV9agyuSo6up95EonpwsXRcWh9bEmrg+gKJbsFtp/qYj2ON8FqR77VKB63Cc3
XAkPD1+IxHM42Go8qRSbekKsFNNR8kgHMf7HFFwkHt5h++GcVUMcfYjnn3O7qwWv
LZmaGgZoZoTdQx7M2IWQQmnydJTa9t1IR5x3M/iz3nhiJItxPqvmCo+sRQM+Ep2x
dWQg6STSuQ+KaXg4Ht2NMk8VpE58QHQ16ndAt67FGpkRrQnwYaytrn6vN+cLebQU
G5EgjwQ/mh5KA7tTrrRTXxJCd5CLI/+IjN8IRfmaG9L5U7RKJYCYo19Y21q/iR6a
8V9IKmPGIGs7v+RXL2G/08oZlFQYoy8XfzhhLo0DaucooDzEZahxkRLQysxiebLt
yaH5Jy2/jPeykPmIYv3hC+MXKIALHfOBi8R6T0W9CyUxx8qRPlFj8zxkbMcOUbZn
SB1/22DbBiLkfjq9d39qgzlkX7GQMD42rr8oyG+GUFz+u4DxVEPNVphOVUvUFUOe
rQca0ZOLmzK4bFEKe5I9rUjivtRpcquLtBJ3veMSn4prk2WOphUE9jxxoQDJSOZ+
CrefOCIz1ArWk2/jUeKTEYb6L3lq/CfmzVZYmvHH1LxSsSgwp8PLKUfUyns79IIx
c4AkODPiej7e7t6N/nWNnJgLpkzlMxFqt+C/ynB7RR0eI9mdUo+flsimdVKApGnN
+7Op49VjWkk4SbTHks5sWHFUumarxniTPV3AzBMwCdFgqKzDv5CKnMsYTZzL3e96
QIhuwGOTXOrpWjF+psUDB9l93xu7mdsOB85+Gwsk3vcHv46HkVMZFow/9mdDUq3L
hPiQqaak4O1sdYdIuLPlR46NZz6Ewd7/SFiu0FzXp1bEmSuxuBXFveiv/nIz3cIg
9/va75UqdmihfAcr0JwLpvWjgoF22PKi5hdFZLiLW08EdJpja19sMmz0lg78LFqa
od6WV9bOzcN/I+TM9u1VJHoGwUNPZwMe2dBfZ/fqWksQ4tmvaxp0JhUwrJpdrNz2
UBc7wwIeaynPD02+yfD8qvTccsbgtEMrOvwcfh6Ui0VzuCdeHP8IBEDdL7fk/xOj
1KmIeodgHBRRs9++4o4NY+fciG3rHGTWRwGosq4gc76cKNsYsDBP1CYTJWQ0t/R8
in3CxsqY5F9fOPi7oikV6++Dzu8Ta2Cr4FLC0wIFQ654rOtkYRAcZmFwvwx45W4f
HVuh/vqLqSpsC47ZlRKjDfq4qm3Yl1RPMtoPpDwc9F2Lk9KFt5kFx0M1kwP8A9X3
XLQcgfKHeO8/lqPy6KODFbh6Hs7lOvv369GOvYkMVopHAkZiMCjUQ+oJ2ZtPaLDQ
lcz+uPH4KyczEs1YbCaQIE3i+Y+4f5x4QPMHB9M2B70mN3UfSA2BS5+y0Jy3w0g3
2ClKMu0yOZ+5CYg/CggDXkGdmqfjqtkL4400b2qck1IcG6R7o+RAipkDQeusDw+o
aGbEZ7QSy3I6CEGHowi7LIShkfU3iZRfmkS953txPd1WPjkm9aupMFjE3uWy4lIl
dCaRfa7sHhpWkJ6HuVpUxuWuzFoMKyAY/Uv54Q1t2VYDeamFMCNV2VPkhtp3m5po
jK+X/bitAV78rq8piHyQo0Cx2cP5LDQUgw3YKxUhEvHN/ZzQaEe62MeBsCSAinyJ
Bmh5NgR+DyJMA5nv5ZecUjfgKPJ/tzKtowMjCovEgH7DE4YUjy4dlLCDp6l3VB1Z
Hq+/CYlUesmfKgkImwdBfejCqXHNCpCaAFlzv6YWBpacX1snf3htUzjq990qF8e8
eIGoegZWCKqQ5q5GWS60i1rOcVwuQHRwUCImJWFY1FBGUqZt6HcRh7ah2CYo1uh4
S7uDJuOF3gNSSppxu6ZAWLAJzdsk3TVnz9Kohr10f5GFgao93e+9ldW5BE8rauAX
uBuvMgTkZrffDvmWbr5l3vv9p0Qsv21GscKX6bn4jlDT0AiWXEWUOdofrGxtjCvb
Edr7BneacD+m5i+rkj7s2UlHsJH3JI2oUjQjRpwFGP1HlMep3nuQTShaNw4XWzPB
c93jKid++94HvO9/0CD5HOz1aH1hxGhjCiWhxGmRCgaciyrFiz7xRRZQPG8RYWvZ
r+67PFUkaLOsCl+yAr3iJI4qdhoBYKnWBceDwBSRSZ/7zJgojyYx/BH7y5PEoGyf
gCHAGvuIjCzYbPAuGg+XtDPA2RhBLlMT4vlO5SUeiNVcY/xLtDs7L/T9cUGD4b8w
ZiqPPvY88x35BMTU3hmP7Xh7TthtxLYqK7kKDPpppkXALaTtOjOcHZ7x5tLHmJtV
d8Jne80QSFY6indFVxd4tMa3Asjqr3gqnycRNDixZNQUyJwVS1Fjo/TmEND/bMYN
r/KYl7E/7bwNG0pzbFAOu3jLxIYV/FCkfUNdIEy+KfcFDkSj6BpSk+rHOnStte6y
W4eOnkDFSnRkOooswsS29HzoPJBLcORgYGQCZRBJP6utEm4Wvh/CQuBy8w7Lu8uW
eQX8+OMC5gaXDuX1LFMBvmSLeo7yZ2Qj9SsLFl3wIsrnNO1ZGt4snLeu4VMuIrU8
pM4SOnjbPdU9RsZxB6xDmY1ECegqT6IsRhRNk9eoAVc6vKmUDj+SY75v8cxV+6fC
+hsIr5LPG05Y230+JuNJmia0MqJbl9c8cqFq+TdVGu6o2zTYkpSi8xwQsJtyTUO6
efJU/uDBmo4L3/79M7D4MiTJkBW09j9UNVj3TZhOlwwzrdMFHzdxQGb2JmMVqqPQ
vqp5V7tihJL8aJHnxhHyU0I4QNc5K+AvWmh8Sk3AslC8t5TCu1oPpChT6V8Ov0qA
ThY0NkCUrtQNsWzqbpKj7OjPBoIzNvcImJcohC8LChWKT3PnbZTEXxvti3HYiFl1
qe6tqjSYTsDxbzJg2CsA/y8gRGbsmZkyJEDkKneECv36h9ttINfqGR2buC1xVqC6
LsP8v9nJVb0nTqCHdMjIG6/rHR8IGseFRHyLFKgZjx5tkCSgAp661lv5inykIQ/r
faV04WROcLjPL4F3Pz0f4CaAnly7Tyl/TPWpdIoOhEByXtrwkXhilc2quaKYjR/o
PA7gCbDIxvh171+1DHT7GRPHBA5N9FyJNi/yJBxfUPZCzNMvS/2l8iLzYJFGUqFk
3qeNDlXZlXRziZP3pkpfSSMQAvbHDvbbLzQfSoOY5392jtQw8lJBhny6l1PcW04o
oGBePDIGqIWneAbcmCdBbECynWnuj2jNtR89WPVL+ieRCqccQqGnQVxdkhCaqvt1
Ek5ZbLZQDxMw26/Qu6Evy5WxIpUTeqT8WrxzsON0nxebja1JcBCkDbdolTK43kVn
gRnkW9ZdTZGKuFwX6pEt7Q//cCv2CrJciapduLR3GJ/NBk8OYAPftqGypG/vvfy1
/TFaxILiGjFdHoTmvuBRya/uemcwMc2wt2WoBd0BentedOBFESKg9uRGDT1XIf88
GsNImZNbRTzbWS5Re52CLA==

`pragma protect end_protected
endmodule



module SB_RAM1024x4NR (RDATA, RCLKN, RCLKE, RE, RADDR, WCLK, WCLKE, WE, WADDR, WDATA);
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Lattice Semiconductor Corporation"
`pragma protect author_info="Lattice Semiconductor Corporation"
`pragma protect encrypt_agent="Radiant encrypt_hdl"
`pragma protect encrypt_agent_info="Radiant encrypt_hdl Version 1.0"

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP15_1"
`pragma protect key_method="rsa"
`pragma protect key_block
qjwx3o8ah6C2Q0UxA9Ejvsy56Xs61Sh4ro56kx1ytSF9d1OSj2rImdcBdAr254+0
4KbrzdoqE1CFIig76s/B8qVkTODh/Lfbn4xjzcB1ddxX1fMEh+SfZueZRth3p67o
wc+O5gp0G5AcZDdHjQ9uLLBIv+ox3mgN0Ukggclrix5mRvzaLxSAt2VxVrh5RFSs
pjbp7fwo2NWgxQr40CMiVruvHMerHafZAHZwG1cFkINvEQ/FgY9Ma5naajpIYO1b
wnKeWWXoxUG/+qCN7wvvGaPSf4kGVdBEBC6WBA8s0hMl7GrBOmwNb4HPepyK2/LE
zmFGY1iK3GH0pq9oNeURKw==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
pgJc+csYqKhb4BLpveEw2VMRWYxjJytvTHsORWD1Xp9Td59O0lMSUgMzFf24Hx18
XtmP9ZbJh9aLOZQ2RcqQ+7c0flRiSO6rUxiRgjJbJWeFK+rTrtol07/NjZd1nn+8
vaCTdW3om6QzzVUARrDfMu9BoOZEAo/zZwNN6uuuTNsFRMKYdZ472OaOWBjtX0kW
DurCqj9pMO/PQRg6gYkwf7ogXghNvV82fxgXSeSwIqqrkj1SrasNY7oAAiCcK5sh
Z7ZreyUxrGIR8JQ0NPzvIWsO0A1PIc88QU0Zk7h1XlhaVMK7r4exmsc3EnFn91hx
JWnK8aIOhZMqlTGxrL/dTQ==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-2"
`pragma protect key_method="rsa"
`pragma protect key_block
W3hXXiwFL3jtT05k5jHTNwyTXZ3v1JhXgl2kPfqQNCwkXNXsShBsEjWZ+VMS65Ol
oVBYlobyxDme7ccv91baUJ9iiNAOy6Tx2i502OrJHcsbsSKmYJkHRcLrvQX5NoFW
cChVt9hy+a8QVqVIvQ78dobTe4T707TZ8EgHwIMO/DXH1rIQGKxM334OFKb9Z4kw
IVplFI1mqMpdtTbndyjwDO2QOiYzEWmu/X0+R0HfbSaGe9aO5hPRd2hGGeF/Hz8a
HUSmucW7FrPTKAtq8lr48XUC3gvVsjDC92abqmvHPHr97bmt38YQQEdXU+jKiECP
HiTjzZyPXf4iTJiIi4ip2w==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=128)
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect key_block
fdlU1jcEq7/SecJfeohmkHvJMzUqEs2eKsDWpMUbF6zVEmwcOACbPt8eg7HWkS1e
AEXR9GEVFtYbSgxFpgFgOAyiZ/Fx0R7Rlfd9r5d7jrbSHCHLhKrWadWp4Xm2YRgy
g2cbmZqAr6d+RPSrU3EJhZ51SUVxo33Ld/qLKgPLN28=

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Aldec"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect key_method="rsa"
`pragma protect key_block
gStpuGD35qrrWzaoUdMM/+jUXCZvFO86nRCowr4xLEqFp2TQTm6TvzpmqXeTxjsw
v4zW3niqMqtVb+kqSbntjNRsUma+F79+VgsUHmZ418iRBeVz7CC884HiIPA/JKOb
ZwY0ySUdBxlRXw/DVBwwik1txlSjiGLQXTeORruLtjzVIMLJqWCUZdkjWU16vpEJ
/CznFFu9grbICG9eom7XB+suaA0c7YveqsM5txyEA4WJZS67vJUqLIHFsaI0VYkW
MfPyCCJncTs2bZlaOWCc96w7QQUSOVDBUxBK3U5vnZxiycxqwMe53lMDga91FYrn
RRbJihRXZnO+SEVx5A5FHA==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect key_method="rsa"
`pragma protect key_block
dmx9d2Int+LHdLAmAeFjXAH49D+HlaD99V+kVv+3efkB05H+prJzPeh8F7EGcPED
GyOyIb0ocDxyqFJjcRd9z90Mk6/0DmF00dY3fOuFRKKBXZd5a+c9zpAJjxqil3R+
3BmWXoPanrV/83KkZDzA5JJQHHzS2BIHpE69YZ4oc1lVaHwvG7GGZyZ+k7pRqERB
Sbm36FIQS3sKH8t0H+GEnLDPEXtIyh+0lQyO+uH9hPBfMApJufrYgX1YUlCeyyF3
wB8PIAZoRRFvO5HmrC1j+z9SkekF+j3qiYzOd9hekeJyWv7Tcrkru2JinVT/y8bz
IZb3D03CuiYPWworMTlXHA==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Lattice Semiconductor"
`pragma protect key_keyname="LSCC_RADIANT_1"
`pragma protect key_method="rsa"
`pragma protect key_block
UCpabZnpOwYn2uhz3In0E0pP21XcnFM1Btz7fukarzQHVlzzHN1kICSkayeJxtJu
g8YEvYwXiD3GlkbOpHZZUOs0l89VBduJwcU4bFPlAFFeC3QCAkm0rptG5u/RN+ak
CsrzzfSzJahmfWkVdaT8GzMLBNmDJN7M9CVktyNOzZ9EkIxSqDQ1cDh7BQq2ywxb
y++3cUII9F1iu1+8859CFarn5qhCptej9ALVHYUmVO8o305fVCGUwbsumGwsjTuH
EMlugPBCoNQONsnsyLt4yGqfpEJP7aBaOYsTXdfbdrVFiqLwGWK+4vUfqcIflL4Z
x50IdPYJu92kwUCQ3f0Iug==

`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype="base64", line_length=64, bytes=3952)
`pragma protect data_block
LfizGAEpl6uj8O0/TT/MN1dlVuGhmOP0Avsdvk/rq0cEqnhsB31RA4nl6wne45R4
RdRLTACnrkhG95+KWESce2QMNnXpUaF93ibyPZCGKt39eMIZqDFAsb7kzsReT5LS
axcUTnAigBrNaN6mhBwg6bZjkgpMt6sFeHW0KijIsjJPqS6bYbJFCyb09b66UUdc
6NATgVoU1Id04ALrjWZ3NZMPS1RI7SWtXzVEtrtT/ELGt5xNkEZLYfCK96vsiDPG
9Dq4rJRZ/d5M9E/Lly3vp90l77QJqKWS6fM5CO4XzLf+5TtnEcwQOv1CVw7zh2j3
PTTLJ3XPNSkRAEVLFWRdYPkVFpmyUt/wELP6ht8gvhMTGt+8iDXaertP+3s8XaWY
PkC9yHq2yY5tjURhgp/TssuwMjhJaOziGVsRiVYXsiwsVcOb34HoZUg2V9qRfWMl
FBI5VZC5K0ULwbZIXsrpVkyJzuSgzW25n57nVd3S7NDT9F+ICWCUa1+SIrJ8YNmP
fdA45vFzstxwTM26U5F5+4+yn8WEbN6qTBGi0wInUni9fIPJivKL63dbCfbAKal8
mYPjUXGTOiEb5La3XzHmOMCmW6nhXNbueRTeBosfUowFph0IH8SeBylIVzDJNSkg
sHaPJGX0iCgMIK05ZBurM/+tXthiVt69CqNNq7q6e7JUmygXPsNu1K97O4GljCeq
SeF13LM+MnRQDdzaeOrcBuLU6cRy1yjo8N2mz7Lf6Ykp8yNbBY4RpHQB+KB9HF3O
m/eKR5ga3VoBd/EYTuTGn5hwjKrk+cfV4nGvHVwhMH2RaxEwpM8Z7NqRfBdywIWB
OxVi043EAGBFDSEr1EfnTiC6+A9eE1DP2cxXgBK/oSeUh3D+hbRANG5x2jXzbBu4
6oaPz/dYosvLxKeal3rLvfD97JbAVuYqYtg7KXrIjO5DSVK6HeEvKpfZlwfv+zWd
h6weImwjbEBKOd5J+vD0Q0NCUDh4GCf/GPs+8RgZWT3+2MbkxrK2tQ5U0zBSNfiD
NPqxFsB1hFOZYJZCPA12eSqDA4Rdrb9RkMufh1UZAPOQjk1dg/2PF21N0VlrqjIi
3unmNEXEW2J8yZavonILPVpJGYv1SndGZ5r2ecDPrLwKokT7eGprDjOG7lP9Pv59
pmy1Nyl4LmxOFuPeii3sbubmCwkCuiFCjyrHtenCP0J9crIqiNXN7zBX3q8tWfPq
+qgqKeJIE3Tudx0i/X8jeZ06YQsqTNUUUSH/rkcufnUMh2iO//pSAq+4DPM7aWTX
3b157cHu8fDoq7fEpWjuZh/FWUw3niluRoyrNDLcmUgwNiRcBWLQ5Xvd7rH3nDZL
m3p6aEswk84fDbFt9EKaHuZb6sZPakTh6T+1jKlhrAMDoOUUWE9PY3PEQ9PT76ZZ
RVNspQSHLzj6Aq12SuoMU9PhfzxVQyPF0fOo9/qZSbY0Ww11FOGyg3QvvJyQpCWp
7Jx8tiDMUUiJQRUajpH3sgyi5gCB3B+kMvkLQAukBQKETHFHeBkZf2L5wksl0ZKX
zqDn+XPwLgyugncTB2ArZ7g4p6ruDR83as4YRxPNMHR9a4CUh6G8zpjFnO1Id3Ip
AXiFva/d24+LhZ/SCFbyJR+1XURJ5aP5kBjTSaMZ6YS4fmo6Fbz8UfcuMcBpeoz5
qKmq71Xqae4MNAxcofeEuvey68/G0V8TIM8HTUohUD8ZvKRp5uMsRg30QnM1ZGqz
a6HTX3h7JxJ7ipdYMzZyu1MEl91xSiozrRJqAep1HY7uF8D9WkYEyauqBevlIrQD
1PrAk1S/KUSv/U/9RRbr81Jl3bFclWEbqpgVGFev00VOKtrIw3vJcRhiTvzeRAH8
k+/kfp9a+Yf0l/kWx5sxhaXzamwHHe+Pwph8+S4M9c5VsfMTkTyyvnyNg0JoOb3y
R9+5PirwiIr4gTO1OOMMF90ZBEM5JLxi0DqLCus7yWGm4w7tB4N8yw2NNE2tObcc
hP1lfyiImSA0PmmMPRfBQt+rSX9c8mggEKPXwgRtjGbiOYvW8VLgfWI+cYeBupne
muEJY/guCeDedono+i17EQmjJLRh7OGPCsBjttMexOrJRHaWDMuMTj2MRbFeVi8k
n8w2X/15dxbxCw3JWZ62mWA2VfxtVV6rHeO5Y6uaH9LKiD+fpynZgreB9I708jsJ
w00U4SaV5qYt25cj2l+u4Z8OdU40GY/8XjsAf+q8K26fKMknowLSzfMe59L5GKBO
SnsJfxzd/1BNk2s+Gf9iOnqodKsAdH6bitwVs7wkOMECrt/9sb5lZ/bn/uWRlluP
LFTVyT5D1vUpF3aBZ0dyxZA//mt9dzNxo7JBD7nEjubhzAtsI/sYc/GMNCINPQv5
ZdTLGD3oWjtC1Z7nySSiodmflnItTG1LQ6hImJwXbR443g+QvDc2zY0F14tVxDR+
vQx5lW9kezIi6JESb9q5wbuXs0LG4WphM+ocABrWCCPgb1JB+wD7V1rKP5fY7SxD
ERyuc7D4/4tsMiWIcIzrug0sKdRNfxXKAhZ82Zbbvwc7tBJlI3xeao9XUx+k6yQq
2WOlD5twV7+awWeTANBJsGOoaw5RObd9CwdL5wHlVGr4atjm73VFnM3QpyuW9Bsi
CZwQf9MdK3nkEpX2/JBdrYr6ivokaRjVPiP2su22BIEnpRSzeZaCRwXKizaAPRpf
PzyLVY3YqBPcyfAMhvRw7W/KRz7xWtDq/LTnPy4KR2woVJQf4973ZoaytssyLKjq
Ou+NvW6l2TUzZWr2YvfrTVUECsjUoFr6eK1J7pUnSsAubD3nT7y3yjMGl1TbsooC
P8rGi4aKiQiIjyFDvUZu41SL8qgDHRcEi8A8AHGiqjU/TeRCLcIwUCQviQnJI5KV
zkFzMFAyjwN/B05ZBtaGUEvvirZNyq5YhpOrO4TbNNa2I2+E8AcmWGwBt0Y3GrLY
Rj/wnm7H8i+D06CAmXHNlAXSLghHhZXZa45SMaFjUBKTnNDGT3WLk3fggabI+xU9
YH/jlqo6OULpvbM2ws0vj2oSk5jn3AlUqYcZECjmL+1o9RoradLerGAhlJIbw0Xg
9Fee17z7JNUtdrAdF7EsILIFtuxhe1arhHZTRxwCtc9W2I++woGiQQyc6QVfJvtL
PyBaC9S3pNAPOGQkYKYogxeJ1OlRENO1UHR5IAROpDpuPAhsoSqV6PVLDXz9fiSU
+fIy5Lr/6HNxykiBJFQ02MqNbNyKwr2g/oXF1c1LJfGvsvLOuKXW4mTvtDjJkSvV
LKm439l6F4ANgJQVhIodxUbX4G9M2vkGXlHfFUN8Z0XHkWJbOizS5pogyMuDH3Cu
MI43Kguu5DoBbeGNDdPBo2R2uRrnheaCaSJ8gqf9+i1CVAJQ4nk53zkN/+QvhjPD
wjtAWvRyK4zqXD30wu86LD53I2ohW8Gj3UBkxW7BM1R0nhqvBe38RTcT6dn15lqP
ud0GAI3aIZuKJSdl3aspqJrtk9OctRPFyMAmCcVhvGu99liBUJbNFnYWWZnwpMIL
Ls7S0GUHcwYyH5QT+mAQaRJq9t3KNG92XrOD+ksE0kWggNlAc/2W/fFRo+pddbCV
+5ZOQjlPJa+0jmFb26zpstBtUKMuuQlYh1HXbakUTGZYFXik4dVRzM/KU+5bn2ag
Ayt52yhFbTZ8PDqoRYHLhXwGjLMaeWLQo4vZAS/QQp7zAjOJKCwumAW/nPoGQjBq
hTMsfzhWkVZb+feJeerRtl9gyTYzG8SeN6nnOSXrgl4H2YmFXNYfsSz2M0yjnJPv
QHzAogX8ew16CMVuR+GdHxkZUUSGKVFDiN0/KWAFBh3odg2eqU1kA9VZGE/pNps1
JCZqfWgn+ZFTzxf91XvskMMkk8nVEf1tgeapbRb2wojbCGnbgq138D1hMFxnOWqL
N/BJjryAiqkM28RGQM2lD+4qpeY7cA5DiqF8fbiFFq0FfIEtQRu9DoXH7jhLTiPB
HeJkZf95EKJVj+0jLWaaIj9Kx2VDZNKgLE3MCYonJAjpNr9kqsBzJPwI5oYtkmhM
ygmtS9/ezgGEwrMYtaV9Gzn40O7IdIFHbrkl+iKEhyexhHI1nabGKuMi6s3qJ1FO
JS2AaMup+LSWGBdpLvBqwhsVSwVkRBxDWnOBuVrxWYWcOpKZe1BzHRuJrEdRnRk5
n9BUk9x7F67afnFO8ke4wjEtQsiUlnGgYYa1hNcfGV/UUKCcjrDYkOS+/hS8oIY+
38Y3NcN4CdpatuD7LVRu3a8F5969UioroBLVs1A1IlUajPVI3D3MHwxMQYpzNBWa
6LwS1DrGRuikT0M9UwpM76TD/zVO4MU6Fo9oOsV/YmnP1jR1tStHopO0f7+TkPW/
u/6wIBUVVXTDTYA9UIINs2AJfUWx86EnREWYONjHBqv5z8mjQwKbGBVgg1qrN8oM
idubyiQIGnxTNSEpAPgewpdEpXaCstwZHwdOPPZoSq62BDZrURMslT+kuAJ1toog
9qlkQgXLFVwZBc71b0BeIxYVzyrsYEgmPvRjsuywe2fGeXm2IjwCpwD41YH1ALox
vsyntHCrIkbps6vUHf16J0R1TvnLSwb3htWDwkKppz9zxnxxTI2yv405htNPXN38
pMwodPNaPaR4LhKC8Rx2CWeQvQS3friwoNjZmMmDksyYZJcKUAdYaMiZKLqx7wOc
g5HdFw9Hmh3q5XkdNIR5ujBsos+i+PV4NqPha12Qf6a0+aHyknMyWeCFFuvFHh5i
/vySB51jkjzKQjntPy/80iOKv48SsGymEW+NKOTvNYLMh2jPjv2UpZaGMyugworZ
svgMzBsYAtJGzYqnSUlRUcyMfH857XW3j0T7xfjjrlfvgoiCkEm+zN7fAZnnxQyQ
NwvTg7KgTT3rwnCpKt+CB+INcdE7EN8cT1q0nBymRkwdOEfBoKq4cQkqKfqUK/PP
bWjN9IouKlcMuXV9CBdmGWUCO0//WahSMAeyuZIsOKDVMTnxGfpLMGuBP5cOffZN
XPyBICA0xyymHYIL6Jh+LxSYGSfL5B6RxocpBI9Fuc/k8MGZURvdHDw5Ce4pDL0v
r6TsC9sQFKZuMOXKAhOU2HMXx8TnVwyAjygbn7zvY81eTC7bPSuPv/Vy5wwv0tuj
cuFtm4zy7LfV4KrHYeXaAA0YEG6q2fRA1DtWrLiCfRBbxuEvltkXKx8sEuXN2XLB
XA+SgOSvQNhnBjsyMBvl7iYa5g4AN4qo1CTgvhgrX9KR5FyCbkD37hMe/nbN3pGx
UNbIKJl2zBY3RN+nd3EZzA==

`pragma protect end_protected
endmodule



module SB_RAM1024x4NW (RDATA, RCLK, RCLKE, RE, RADDR, WCLKN, WCLKE, WE, WADDR, WDATA);
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Lattice Semiconductor Corporation"
`pragma protect author_info="Lattice Semiconductor Corporation"
`pragma protect encrypt_agent="Radiant encrypt_hdl"
`pragma protect encrypt_agent_info="Radiant encrypt_hdl Version 1.0"

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP15_1"
`pragma protect key_method="rsa"
`pragma protect key_block
fgWkVNN1zw9SbAmWP+umZnlmoiPsrtk6/8auz9aM8y2zkDInAl6X7PXqvA2Ecmvf
vd0wWm9IwfUAq36nTWG4KgVJcdEaCDykih/eTyfrihM3x8Geb7g9GwTtcKBU4PQY
AWqWTk9XBqRu4dWzgWFbw/j0Er68Tb7F5ZVLwncIxmTcpHXb/BXzF/m3tZ8b9mmg
0ytrT7ALGH6291mZZfr6DHxCqfIjW31fw1NSmZJB0mlrXRiskey+uHq+yCw6PfxT
Iuw+eg1JbqYAPfPWtYVu4VDD5l9fP4pV0FxZL3Af7qHynS0xG7V5wOyQXlXsFyKy
lZb021sFI30kDUJGTtktCw==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
Lw92q3Av1/AzlVc7QsUIUP8GCA8pkDP+1hHRJtIqysjtCCOS1Lo8+WYL8HP2H1h0
QPvfvTMizZv7Xxwo8/KByLpMjHNrLUm2NEl+lx/3iL8u3Mx9G64myEESRgqv2jqm
zRm9pn3GUKELB4w68kriPtRyrurW8AGFKHqfGdJlfPHUtOerYFzFEOR3hh/F8o0T
+463XsTtFTKmgIVoReCPFb9QUclGSR1AzUhQT4x1ohQ9UVyYOGrtw0XmhRXgJSha
mchXo62T40cDCDc3tbwiPb1cccxmUwlsGqSr1AH77Ao5PmzImgswUa57pfGmuc6l
f61uw7pFiiuZPIxpF38T2g==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-2"
`pragma protect key_method="rsa"
`pragma protect key_block
FHl6QlGdyMMjB0IE0lHhzwNMSZpv41hG4jruHrzX70poA5SDLvaXh4hpdmTQr8Zj
8jkcJ85u++W8x/xXiDc2379vtcwr/4J1t7mvTtRtMLiJ3yzzH/drfKV4nQYw61j8
wmR+X219EFo5x14itOHhk2VrWeHvxN0+tZYiQ0zM9levgfq3OjYT8lYgUH6Wd+f6
wFasJFi2irISDrfvFnof6JyBIk+5oPLnlgwP93vEnqLU1ClMvyaPTebrLLnz5RWa
5Ifp+yjZrzZ+ankySOv3EE7sHia0NxX8Jr+nUz1L0F08AZ63s2IT8s1ssj38nXtj
JQrWf+/dhCu6uvMdXMUNrw==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=128)
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect key_block
lFr7HNdaMUNtPRsdSWyrnfAzyT4kYBSre1xbnWe/sr3TGVqFRjQFeLC+DoVhCKXe
2C4LspQLacIsCQY9pKGrBh1+X6wydz5mD/lNp2qoYqSg60fZEYNWLD2a7/8LD7M/
D/4lTa1+Evt856gzLru4ATUrUOKZqfXZqCsJwRTd+CQ=

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Aldec"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect key_method="rsa"
`pragma protect key_block
p7bG1N3cnM5TYxX/dwWAhZ01Hjss8e9pc6BpigQIf2zeNmQ6D0zqH6d3aVNoPAWf
GPvs2pef3OratFLt/HFOIVXnyhUDJSsZWM8BcChcCccVgPjc/Bv+hIORqeBzMH8D
j/nxcNARo7vhfhEdMASia7iwkePHyKfb7IHgKoPkyy3xAj531gfI6t7ClEiTchox
BTPdsoaOFL1i3MmcN5WiaDLClxNiwj6Mmzsvtm9QoCQporXgdcTFOYNjjX2uohuq
kGpXt/TxssKbITEET7HDIO0AapECObLMMTm7Uezt5/cSW1K3K9qfBZSI67zQmo0X
LZti4tHdhBeESHSsu2vOiA==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect key_method="rsa"
`pragma protect key_block
NuJx13OIDNldQdV4CAHrUY+KsU5MUdtZWGthtbGh1Wu5g0jr1zFSVRf7WDUTaFse
FoeS4rhdX+qDeSCzRZ53sF29FrSCbhpzfI2XxuuZRUaobMzgG3ab2x2SS6LQ++ph
ApJ5iS1v7/C+0Z1E94+G6wQccH3D0Ei3fc5znPJm4xIhNXWTG3vcZBAYsnNOVFG9
38xj4PGkVegh9uVl9a1H1urGAGBR2BwcqhSxU06MrJiOTw599i6kwvIp2ZP3gpK9
yFLnLZRND0/ShhKNS0+g6qTpSgZvusitlonXnGVChTulMeyXUs7Q7LDevjUCwstz
mVr5pwXbzGu04zOCK2CjcQ==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Lattice Semiconductor"
`pragma protect key_keyname="LSCC_RADIANT_1"
`pragma protect key_method="rsa"
`pragma protect key_block
McL1qlbUjeUYpHC8Xsfd8gNpAY5oW1rtvbWwFdXZfF6StFMt4hohrf/FwD8Y7/fs
Qd0bmb8bjIOsTBeD3nluCuoo0GhjMTly5f+Z+KXJ6wf+66mlASN2iF9uz9WKJyH8
LZxq1CMheEiLxAgeNLZ43N4U6137x4aMWZ03EV1dILdY6siOZcpfFQ3vq3sLgK3v
KmG9o7pL6JztjGc2L72Kw79dMMSyW0vyLbaBpSrWcM47DUMIZkdGkENDriZqpk4G
E+197sUFYc1WjLwsarw3aBBpcXZWQM9pP/SLyxjFdOE3oRohC6Z2PCdJMJhO+tT2
f+R3cqADMs4CI3/AU+4q5Q==

`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype="base64", line_length=64, bytes=3952)
`pragma protect data_block
r2F7Z2XctzxGt8R0rGMkm68wysGGNb+Oju35PVVO229VjtAPftHvtL8hnrG8+LUV
hJpX0cPpZ/wL6AhxkSWuwQTVFlvmYTdvkQlvTz0Igddiz91EdBlMyNQxBMkxo1wx
21VdWxWa3CyGqoRVCl2IS3AY01iDLh5I1jCYDLrc08EjLxXXu4cZs0rNbOyvBUkB
i0OYNwJYqJElCb3KxQcO8VFP89R23zva7iI7EhQ1gARXJtKdqGZJKYC/IsiEd2kB
yYwcJEUTky5+77FLzDBJOjg1diSqfwRQw5G/+KvoFGWh35nyo1p7+/LQuVyCBd2k
FroJlknkg1exRLEUhPfFEU9BP7B+hxF2HF0y8twkzJzjaFjztmmMA1yrHTMSm6PE
D9b0cRmsmxM8algntTO+W0VG2A2AmQH3Oylb/YwEx6Ud2Bry+oDxAVd19dmlbprb
n7qogQqrvN+/h92RCDoLE9Pq6+kJyl4yjnLIGAXf4+0Bf775uOndzVkVBUCPdiR3
muRoMASk+rXP0eJs9kO+9qDZmeinUCSSiJMFDngysv5xQO71DEEDiQH7m3RLS3xc
RK6e/Nio6Kq2k31eAw21OZxyWwna03GRVqG968vo0g1g2+qjzyir2KU65yHhHzPy
sB4HT2mqdJyrHdEVbBWo0wNS62/ZxpGFvSJjnT05SqY9ZUfDKy7mw4y6rYpmXpNp
TM0u7zMkWqFiUrFDv30/jYlpCRi+uVysWLW6yqKMkThQoQ8CbeSwswE/RaGKmG3Y
fvMDlh3tttYBpQGE+0Xe6f4xfqr+gU2kxnYImX+0ivpGb6QD7fRlkpbsrAURj8HL
T5Xg8onrmldhuTIAv4gtG9tNrwrMa3IYPdE1R89sRd+ncKiWB4LDWhyz4QgzZCcq
AvI6VxTlvypoIS+GkSau/W2eM0sAOz/taH0lBB40II8ua+RU26nCj3smkWpK8z46
PSLZA1B2t5f1+eC8l+dNGCzjnh/DIhVMfd/4GAZQmNtkqEqRS+RiMFPUYHlkc/JC
rGgUKxLOizA5cMpC7icy6Ilwu8fARhPkb6uMpLaEbRMwLsYwZQv8V4wjoaLX/DjC
s3GvsrMrwVsP2mY599V24Mgvj9NFAlLu0Ov+fd+lou/aw4OEALs2i4pRo/6PETQw
9Fl07MjlN/XAC0DxJpj3YTfKGeGzhF6NB5stNua3AoXl/9wQqvJRGLJSya/PERgp
Gt7OsT6ilo/uOiRv4Qv+hqePZeJ5aEM7jLST74CxaMknMBGYP480AuSJqACIfMT0
pUacKRI3Ubw/XpbbTuI9lcrLLGHqy8q/MxxdzXRvy1+T3PcmwS+qZ2twNXkFTKAd
+NanqDtNmeH159a9O2UCYQAR8+ay/5KYdemSgXa7ojjd1uHjyQfwItJTk/Li2yPr
/XVoxkvYcwSJ7ohUcNkb3j7KPOsz3KgbPro+Yq3HpMdIeFAy8KNaNYqerVuq854E
dM8k/KEfJErg5p9GX4S2lHWVpqHTkSLR1OqbJIQkxsWEAIEhsKebVU3UCTp5BZI2
J7XOTdHWHEDbIQnFPCgj4Rw7jJWqKnnBr5oLJRpsivKEdsbgR4sypm9pHLduhR94
wT0Xq4/++3YVhhqMRvnbgWfYssk/RnsfNqBztveIM1c/qwR7JPPlF6uhJF+C+LmL
rINraS5rN9j6mjHRHvbPAB4dK+OUw1gf2p0DknO5psGbI8k8uoX3UrK31mQvAQzK
zwr7LT3iLiljGFjdQKG1GN7v5vsYxsiU7+u7BKwTZajacD/ZgcXhcQ66Cr+Y7Gq8
KGgcY50QdzvcfcZThz/SQVL1n1fXxjlkwj84o7KQRrLQ/2YGiLnuZGNwhXRLBmtb
jMikUbQESpZDvG6sqsAfJEnhJVW+b8mEjxa3CMhqWQNCE2gu/AryxJgEIFsQs0Mi
ZP2yBnwTiT1wUN/2nWHKUiJVXY89EYFpxVuvtwRN7g+u2AGrw4pBCbHFrT2NVWzr
XcOdJGXufFcIsVDr8sg/8Mgg6Cju5hh/JqWWtpcpF/s6fKOYbwQNcZhoufDtWcCy
iJT6XTI7xfV1GQc6omuocap7hZkcdgDY0qmxfOt6wa+IO9O13XpY4rWQE8pLlE+D
cBdn/E0dfatGyrraCr1ND/uWuTQh+Th/FmSJ71d4qK5J2pGMVHKKpXtjCEPPBwao
Cs+s7/MRJOpjbqp+fhEZahpGY79rXWmJ2wpM9G9izWMUgXEGY5nxwsH5Sp0XstM7
IcrztVGYXq5csmER2iRhNYvWXBJLEvyQ8RP/62GQgREcWCGEJ1RBifpqpjftVk/s
wO1FjsP0U9XBRDc2UfjuKAMML9etlB2IMyGfwwMSeNNT9SyLxdpl0oLB/8F6/Qo+
e6rKG4zkEU9cIhNg2hcaeKTwh8KW7tP7nLqCFjGMWLb4jHFbM41k1vl/v6NXZmI+
dPWe3/zCGxv+pKpCuFv/u3v1sRLFp2IJ+N5RjCpuNPhC1JCoeq6qOzbRhUuGcQFJ
ax5FPDU7vZMe+qrJg2CB9xBD13uXDTFl/ColC/Vz2GVrJkyl7ohUPVQydyP1ZKG0
w9sXi9QkebhWRqe7+3JlvYIUkU3Gt5Op7uyUxH4Tc8fuETcQx3s3QBBcVm3LiJ0d
Tc11td301mfuDXeVnSnq0ujTVTqbvygjZIpgoS3rm6J8axHxUSTtuRaM8d5o12kT
l7vNl9yAVRuGYKyQZKTnwg4tzR/3TrlRI1+xFNrIpbJu1e0VHHWOJRWZljeajqxR
D3sUGMQ4HwNxTIJDioCmMCJTA/PNNznrSbpZXcsoBIl0nDE65JT/h3ENsGmgfkfL
NIzlga037jtIjBIP7LYxzy/WGyDq3rac1gZyijWFTztbStd1N11uWkU8PwSh0+9q
elgdOv51pWzM6icTqXMjtW+hFO+fgY/WbvxaXA//9b1Jt/K6OUTUMzuUWcm+fdd9
4hxVMuSQf3ZafrMki3Vm3eZ4Ia6OmcpgoYVDOnmkGnSIm7KSYz1Hm1ExbVcu3EVe
HwcUs3mP/6O/DwzYNXdvAf9Abz2uGgRsVTgIdIAZAjnQkRLrTY737kN/sF6RyxHQ
yJ6/73YAJAaXy4KvGbJu24vJKUViQ2tM1disfGyP98AAOP+ti0LRdR10oAo6+a+8
nFx+M20sxQ9t1QlI96UnoB31vRO5CNJH9EkBvB1ZgtO+hqIMWcgeOTlEkUL1D8WL
J9j6iajDYthg9bxBxDnNdRARFH3aotrqOz+mfTd8Z6Uhb4CQtWqdzvj5RbLuIHAy
rjGVXMMP5GFopaB3dQv1zUrXHbR0rgrm3mEHrb141AtMtYfK7Tgd3uwTemITzWFh
WGRJ4qEkJRTFqmD+HNJ6VMW8s8Pa4DZVYkWs/CO+YvQPyV86qpyvxhFWKJjDd/UM
Fa1aB/+B+vwobo80nWoND/qKMm6Xn8aMffKdEnI36+v+abYdjrf7gToJmaHEcVDZ
GvJOtTKOQeQLfrWqIOEUAXOGGqXZ6YvkqR8VRFFx0s45wLxWSrI4RJWbnkLVKx7K
Gv9YYVQFprSkTynDSoq7Z3mAV9gLTk5RGaWb3ihVsgyUIqzwdIRpMOlykMarzddu
DQFfuFLuQhEqvzINgwRPq/dADuloXtnqRf6Sm+HNwLcT60Fu7Y1X/b6amrOev80Z
up7FhmVoLAYhLJxMNpYkmQGvcprj6KJQF7CpJL8tqhY4e2TCjMAKQNn2crIe3yo4
QTFGLf+lEtu6+fLFy7aWEDrbWkoiF69yH4ZQ8k2LnRXZnXKgmzQDzUhjIZdDh0j9
PlY09S4zZvOmD9cfxbX2TOE0dAyLjS0+B81FYwv+CpmMQPpgHqucbuBuvI8+ldT5
/z/pxxvPJc9HnL0CGBdKs6zLditk9oXKu6s2vA11jnKe1nWrnTP2fnZz1QHJQM04
wNADUsZV0QWFy6xaY6YaCXGrJKJTsuDhbzMWwQDpL2m61ree+HmZ/n967ZL4N5vc
kkAB5/+MEvrt4yAstrXxGEahqy6LBLa3HuRJcGT84rqnGCGk2eGY1lB75rNqqufa
2OfmWCURPZjRfXUogN6EoUg0jbiwmhfK2fNeAeAIPhM91+pdkaOcsZV6ySC/LpY5
gBgUQVIebisupsFcBP/RH0HKjy1JTX4egYQZ5O1NfbhsWleo1Qm7QsxuD2zPjpKO
p5mzZzFRyi/jbv3J2qpIfORYyYVWaL59fg6ayNxTK2FI4h2LKLtXRRYDHHL8ADhM
uwqrajwRglEByGiieESrk5JSeECmwyEkl8G/3ck53/rZXDViDgW032pyEyx9oTgk
cTAieEbhTCj41ot7Y+lIIFqQFoU7sMoxXIet1C69K7O1x+Tbnz65dQyaVYOKwD2K
XwjtuxuN6beEULzIIPrXbUOWPALUgDY2mdE3s5wSpt7fIcX8sjoGQAJycWeze9BZ
+opH0cla2TqnuGHLSIiWl5mfWh//OJe0RUmz1WPcPup+zlKaMVFiXRD7tm9vnF8G
Tk2baf2GtXRgxD8M7piU754cWPVqbiWaLBgIGVF3ddia5kUWd5djF384rm9uorio
b8Ez+cloA+aQZ1n/8B6eyykK0Lz4aZalwGELYjtM10ldr3X3S091kAI478XhIf/d
g0aAw6eHxNQBT2e6ZdxbZZTFfjF5OLH7YuMMbCtgPRKGde9yJZZEAJjpmtaKgSSP
9jKIs/qLLQT7NyiMJYpoC8mZgaFIDfl9lwQjof2xsa21plZa3d15UW8Mm70vrft5
eD6v7MeZ16Cu30Uv/DKU26DEPsG7OC3WPR576fHHpAn89oFmBoB35LQ809roAEB/
Otf2+5fiZrcpRoWtjJeN8a9fZtDz7zSOhNO12CFN+c9lvMx5SGX/CDH/gcbogHXA
QajDyDuhVZLUV6kj4YzycCEypxxY9EQ2WrXiHMT9WJY0rHsH7U+r/EuW3ITVo5ux
TjHhELjhcV/+o/klAiAQcK1zYLsiim3nNaMHFNCLFbPH3YkQQsie5muIuRwqQK61
2eWOaUIa/DJK08N4wE5dKiT896VLHj5SopumJTBU5KCEoNVlW38fvTw79D9cfyWj
S2rmbi1SHxIPZvtYqLMYiSwDJ3uBshNdqfpnQYtnumn25gPE+fpIta89sLYgPKHi
yGYwPJ8CJjA+zqNYTap/POrAOshtWRNdy1WeHNZpJkJRV6Ken3WfNX/MVTZ3AYkY
yjkqjFfRbhkg1h7awn6Fn6vuXBNJ96HkxzsbN/gmZNSSU+yalXhrDbMFPm0qwt+a
OWkTWbRZVLLhIm7fzftELA==

`pragma protect end_protected
endmodule



module SB_RAM1024x4 (RDATA, RCLK, RCLKE, RE, RADDR, WCLK, WCLKE, WE, WADDR, WDATA);
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Lattice Semiconductor Corporation"
`pragma protect author_info="Lattice Semiconductor Corporation"
`pragma protect encrypt_agent="Radiant encrypt_hdl"
`pragma protect encrypt_agent_info="Radiant encrypt_hdl Version 1.0"

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP15_1"
`pragma protect key_method="rsa"
`pragma protect key_block
Fh6HFVj532TZSMyyq3YpR8anELOZ+1SbzzIWf5GU5n4g6C6pPlxoA2UQf++WsUrw
wbZUsZkG0q5E0P5xm5k7aedPmrvhX3BXFCJhTER62+8qHWGxA3HdP8bB0Y7jZumz
Ovz4lfq4GZs/fusYGNHs6WiBu8FxkyE6yL/SWf5cdC9d5ODs4s231dBs7VLhsc5t
Y0lJf7u5nCqhi338uPzxzjT0A7qN0sVFmh7EQqr8Q4tZzNqDlVNY2bjUF/AtAwda
+UcSbN/ndrjkbGl7VE6PlBQOoW2GI8Lb7/4gbQkfE0VesFBxNynM77haQEe8fMXV
Uv5lsQCxAouftYPmJoo43w==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
DXfrqDB3oTK8GMvqNS6nVlLhgJgq1m8MTFyBSAgAtX0vRuvuy6Z7nbbY8HY/3dmx
0gBC5z9jXILPnFQqSPW5Dq8y4Ho38En8Je4dKxIze1Mc3kLUQkaA1ObE8F/2sNN8
k4Y6f+CEMYDX4VTwr6a2K5jFclOKjz7kzqynXnqz4+Sx4skSQezKaCfTfsWpQwHT
f0QA5vmD72I78pl1Mkkl4Aao0QAOHhOqH9L3LWXPJB9fHcA2dvhYK3IMSPeqkQDW
StRqCmcHRF8zunk9o3O/8+KiCx1rchpsDn96mul63Ye8U6ikAxTN8m8Djzs3Vzvu
fYstopC8zGQQ5zMs25ETpw==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-2"
`pragma protect key_method="rsa"
`pragma protect key_block
PQwPlvchcnjlLvk7eKwVHwBPVzBZXGnAxZ0EUfFC53pnAdVvy7WBDgisoNzlgMdg
U6gZxPTzrvGiOGPEKJh+/BY7DLIoA7bg7TTEnQN+WmX0UmAXvIdhtawzg5PuY36r
yeKrGF7tL7/SP//GLVwHkiaYeQtqJoLtx/jfnuH2u4qlKrt5dWXG/S9e/yyVADZs
KhzylBv2tgnc04hgCnWH6UhQLLRn5D5zU/Sy0nEvkS62tkGp38zCaUCqwaCFUb40
Zc9ZR+hgE+tqzdNeGW3xWdbC6EUWKKBFXiSJCIV+WFNgKDmZIIz4sg7jsNpi5GJA
BLhdGv/xXowZ/+fxkwk0lQ==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=128)
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect key_block
DYnE/adNyzl/MJPavtq9xeVSYOvFe9NqTPDV4/j3uHkgq9kdejOS9G40gew7aqwd
FFLPpicGgqI1SgRSy+AUsDhM0dJ2DkPezj15R+zBkwMCkWybC+Bj/JTKu82zPd/2
R6BeNppti9FAzXizkjnHA42jbR8ET020GmuPyQtr6/w=

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Aldec"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect key_method="rsa"
`pragma protect key_block
n3tWdLXtck9tLqB8iHQdUvvR/TdJVQ1ssm4E5tl4dD0hSE4FMVCzd0E/nRtZf8Fh
k1jFBqVjmRbzRJ7geIU04UOw5AEUn7dz6HziOUg/qJNYDYyDj4DQ+7qIERkIUgPy
kfsMcguNm33i2o0q/MGNIq3gmthKslamnBL8ycSoDGj1meZFMC3TcyA7WeNBTfVo
E7OsA6ZejGI4EdZ7qK6b+Q+o2OvvPJBdcQO+gKxuuGUuk4V21Ezxlzj+g+UiXhIn
CukRYa/b2KtYrH6aCtjCBo5f625Hieiq4xSLzUcDKTLNd/aryrVTgPztFRxzUqis
4uY/V2K/VR9gXlffs/wFSQ==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect key_method="rsa"
`pragma protect key_block
aIiVQTgcJWe1qaXecdH23ZLrcuc+8jmbbKG4cSt86DMpyAOz5Z79y3zdfm8wEgxW
Nh8kssWZQWqd0+tV+ZyCU7h4Bu6TOf1hD+UKI59j2PwteOC+vuXT4sbNisiDIoqj
ncTOmUJYJRMaZYVNbdNlwIT2wPppNi9UVYaW3c6c5Hzy17AenbHNIfaLh49R/JZx
dK4JB5GpyQ7bd6Tn1BnR57SfiXM3/jSNYs0oXpMe2nMKumqVyl0jXn2TpVt8X4km
sD3tvtjv/1DrljCK2xD2oQiv2zbSZgk9TbzjzNKpQ4z5yjto6Nb3oVJzYDYo6WU6
+FEPlJLxXRqkWltIu1ny4A==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Lattice Semiconductor"
`pragma protect key_keyname="LSCC_RADIANT_1"
`pragma protect key_method="rsa"
`pragma protect key_block
TpfRhlESwTnCa895ZXBiMA6DPmggNgY6vBN8tQNXrSHNFWiRe7cqnJ1HLjbquXD/
GIDgYU3INBajJUIIZZMyv8SqK24I8r44oQT7/PVxQQ34bzBIw+BR9cwJPuVE2l90
Bc4r7nmsAfhev+3M7IC+P94HnUKupdel/rCaPyxs5vZd+q3mCbJx+WtRf70TW/MH
ICzof2TsitWzpWltXIfQCmaAvUE7rrdjLkbRBbcSiRcajehEIREqXJBUU53qA9Hl
nzkIwxHtlFU381Os7NTkM6z+WN3Py/MxBL6VyWmGv1H4KwLS9tgVhy5P9hGJAW+9
fnTE9ja84Nitc4ZWlkyPyg==

`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype="base64", line_length=64, bytes=3904)
`pragma protect data_block
KUC9cTTaOSf4aZw916M4lPfB8SHUqolERTtO0p2z3S82i5EbQRtt3aCxkeTyjhzL
5UL+gOLIwKx1BOd1GdZYCk/38G++xu/SrCFkzqkYB1+pz88HZqPOLFvmp7Wqo/59
J6QLmyLUa3d7Sl6oJM9s6dXVrpmVwok6Z+Jo2iXWLC5tPZjQovHmonv03sP+/cT2
zD7/4yf/bFrtoTLnyb1nA4gDOagSXqgnWElq7UzpkC6/JLd436fqSQFoyFM02kaK
M1GkJmuk3s5GNPLcwuEaQlK00wmPWuY8lDtZNsWHyDgC4HKNH6m/G1/bEiCKKyxy
iLZ+hCsSk/HNdg7gh2EGSOMYfqTKNJbWPgWSOQKUo5E88TbZX5q3gkKi/IRvyu5P
Vv0fOP1dOvBuy4twU0VzpM87lS9KZY3vI7l3wmqqY0TnpMp0SnX8XHgYDRauhxzm
gXMid14HD7ulsk6DB9xWoLmXiv6b9On32DActdvg1nDYWwPy82vd45M2kGfWePlE
Wi5bzBLX/CBfzBjdEGl6H5u/FcCq8Pw1j5DpUijXNkyKDZ7lzD7t9mLJ1GSvN6Vq
8Buf9G1zytQ+Y1J6yP7UJ+1cVO08Apv26m2rmMZJ9irueiilb9yU3CzMHPUmr4Qi
aOxSAmW2jNnknDlQIGv07irShZ3f2ehtE2kL0gTI6dTpWBJ/+OJ+JVtf6Qw/PVLE
Z+Cw6KgtCbaUYnYJLy67s7vK5BrQhmkSqzrslrXUB3VqVJeJK/H/TDR6VxrzEWWV
WMtCar2DtQbi+lNVhqA0OYDbO6h/yqUzAvMT6+FAkHsnq+BABZ3iVwHER7Iyr7SB
NtKg/W0gqSeY+3qM6oarJr2eYDc/uBxedhX2GHxnce4dahY1QHw+MS5Og0P9TXxi
QcELDP2Lw+QUtU8XxJtA75hNEzultc6zLHHkRO6GwOkn8w9nO7MEF5ZMJOcOrqDs
y4WLKoPXgwDqE9/SfrZSJ6Vsv8ext0CvRIbSHFkd3gxYsA1B30DY5WXJBDKptOEW
YWwRlmVKm36KVQMRAzCoesTGxR5Q0RB3UeEZ03RomfN0dXRCNff8IPkWI9CWw7tD
iWo248mytHLT/xn2ir8LuIJq4eamMDnwy0iIGK8q9XvWKhxEBbAFr4Zy4RtuhG/v
ZnfLYPtXsLGejIWutMr+0K3FZmyy/wDuxI7owl3Vb8BfS0bzN7zIm/Fgch3cEBIE
JBO+rDG62ryMsg/nYYBg2o0uH5q4RxyzdUjUxnIXb0x2dIBd+aOmdE1xUBI62g9L
93MEsUvpARbyIVmYM5QHyvrPrzPBjjQOKysQqqZkFP0nhZtWrmhTmj7gK9iXK+nH
+/Q05juUJ8iyHA4x4+MAddsZRUgifTvIysjzNBOSsJnFQFOEKfqM8fPa9JV8g6WL
ExeOSxZaqxv+AGDuaGkoDYSkA7/QnG9CoHqhzjj3AEkzOzCRK7jOsev3+v/+TFbM
nN70LaLCXN3ohCTO9wck+ZtqtuTJvghQnm5vp3dYcKvwHdNDpN7RyApB1cnaLj2r
3VTQi7kSImKyfGtz7qSm6bZjv8Op04qgMYVzNJjL9L3sDX7MC7D5tgHj6X5u/Hzj
oy54yQlA7gBH59fczqBcj+68ypflnQV0IH5e4MxRF8dW/OOsJAN0jWcoJQGdXdvN
LPkxS/kARDeRHFF9pYSUN06RDiO+a9zgSF5xopTYACYzb9VC/6JQLd76IqnB9qXQ
hPlqyNHJoDF5opinlVcFwkPwf8m0e8VSeiTyVBYuRp5ds6M0dprGhQsWxd9aHxfH
zsykHJXKeaj7mZEcwMyWPVDTWHh4H5mYQceFa5Df3ragoCgTk6KOO/BOue9fsC6l
XzfDQx/BbHwnUq3t4tfGDADZ5pDplVAb4x+62IIfkV/TMiQiMI3W8AGVFGa4x4lW
Var+r0nlbcvv2QdvsFLTOrAMrcbK2B9PpefTCkbteBJ4L56AoSK83cygg7Og37NI
J/gUdEMz2o4lgqPJU/cmHQN2Kg/aW6DPY5TGHCsALHvNMb72g5S2L6WIu0cmi5Vy
Z8gxhzSDJ/XlTE37AafrXha7cjaKKqiegDSfcIcblE+dms97oB3XmEoRk3oEKFAM
zUUj1rN/lFQWNDYvlinf4rs2r5gN1cxAxLT6x1/zGA4xpzXLx/F+T6nwnoj0DDa2
lCqOCe6KpV+C33VacFETBhYGHlY+/sfuWP1iCBKmwMZRUOVtVb5TNO4EjSQV1Mti
coPD8LC6kOg0AMIBRVyiGHcCDdtViuywdk9W+KucgHWtgARsvHvBkNgXg5N8A/5o
9UsWHvViWSjccU6UxlJykKmq3YtorWyCG8E7oilcdCSNSaRCgiWr1T+ONZvIm/Cu
O3E3elVjEY732oxZ7tjCxKLg7fWKaBXEGXCUoLeLFZ/iWun2RGixtCNkvqKTTyx1
IDPErehfL+DEDdu1iXte+9I2XhRNsI5DwWySWQwf77jW/1z5aWs1bBAS3c0NMMkE
1G5LWtQP6wcCTe4BAa/Lo/oF+XYfWTlh1RyKfiM27rwaYB6x7YY/qpdnbDaZEMsk
4rQMY3SoLrSKRuK0uL7QfwS7xCU8Ifhu6TA5WhA2ofVzktT9axnL6VcWu/zttLzk
JNQQk6thsZVJBivEnu8Y9cg2/JwPZgesabRiEi//wUC++/rzWoAV1jx54E8Kd/Hc
A/6a733rOPnZ1Hnt1qKYQ1krn6OwAVWEtiHE+Vj4OMi5cDB4M5Kle6wQZ6bwAmgC
ngishZhorWD20cslqwb4R3xm8QDIkqzSvyweQ0e+3R34VFGiJK2n+thyP0xU9PUE
6UUue2A7DdErrQAm4amrTE+6ezbPeZWi5ix/lfGjm6a79wdwo1mhtKg0o+q3v/r2
Kz/9gqqXpWmrKl3C4dkPwBGB22wFrm+vdiIhO5p4y78BCnnKPpiXUZ2P6DQcAwQ6
yzX2++HOJkRp4Qj+97xiXii3IB8J4wJ6mn3fJsQPotr0YUKOcd1FQ4arKBrPEax+
L4Kc+rFQG+L2lilVXAOgY2Y6D260MdYT5WwtKxQmYAPgQEb6+mL7YTOMqRkDhEIC
eEDCqYqC54HCj2kodW9qIU5zzKYssP8G4AthIvLsF4LaO7Ie+Ny1cAwB0n3pzAQv
BUlRYJDB2OXmiHWJFdccPQDpiGKj4qFEM8LgJZ5bKgKg89fhJLdmSSe4Z0BEbDnt
PcbzmdyoEbiutBf4kBVcE3dMBIFAGFHtCxbj6Zp6uPMJGOD8j2NzxG/dMzLJ405U
690PrEzHAdYZNW70LV51WiklFQYPUd09MYgMYazeR5OwVkkjeUhB++RQddddoMjD
KtiwMiqMLTRedDoGmTpOuF2MTocWgQXkC7p/VzYrrm+xx7/rJ42X4HNPHjckN9bP
JKSd4cgwSIk9l9p1jLIFlJgYMwdj1C7Fh48pbA1zP4S/kAF+lGjeOQb52rCVhBWQ
KhnqeLU9diu6+ZOEdiW8w1WGY05joh2vIOBJRm5/uJN/EUMgyc/mcqr7U07p2QNh
pZrCvttVbb9fyiRcpqTZt2000nbLT+lqYWuENjI+0qGLCN+UddgWVXr3m44zGouY
fB46okwxZdkQ3u5b/6Rf8LGFdlmYhuVkoObw9zCQqb0h58oABSAm4isYP5+echWn
ooPgwn603Uum9WOjWojjoUoeHwxlShAfq4QuyD7BVWm75rJ5Qw5rf8ifp65jb85E
xfjjskOsVPy6lmuBjkaWBqrlM8C50+pzl8NbyuBEf4XFOZtbJ7CYR5MGN08jKyyq
qbg3NM6z6CQHjtlIBLOVLNx8D/3RmAgcRCutN+3O75QFSdkGfWZEfZHAXiw+OHwT
hZRRPR93fGaS9WcohT+DxOMZ3COfajFJZcDvzvsujnv80LBpSDXZwn91JU34SV6N
cjphVWxEIqI2qjxxXr4jEoRgSMN/xINRmlS137J8Y7siqpsX2OJBhhAhmzdTOdi0
rvBVkk0xhHsN1S2OU5AvJfIfAM/3PmrxsMU+lb2s0jFtnEji1RHDK7e0Buz54zIf
ygPwUOmNBAJnEN6nggXK/LtzhAhpr8UAC57HipFlA7HgvHa6jbV0Nmifq7jhL/Yx
V0qu9vQcNffPocbqZeuScWqJ+1jCXQ0X9Ykh4mkEtAEVrjzMPiC/oPzZ18B/V9XM
TY0+ubxO7fdmf2K/G/TKtNVboSao09ZktsXZaEwN6whpt6MkjmjTTxpsuWjDiLQs
ynasSSt7Kl6SrPbC589+tqY7jaUU6T/ZyWN6ChSXt2KoA3c1OBosVv3gZdvhDljl
KONYZMawrxfiA1GPd/E1LvlPqbl2P41A09aXXD+Pm6H52SsYeXlWn/RsjR19X3Uw
NFPihnFcRJ+InVDmlFA/r0uAwHYFY6A+pCgmFY+Cw50LTy1NCRmLOYcBU84QtQf+
IMpeqDaiyr9tRG6SXzPlm2yt7/tLmlNdw/05bZAp4K3xj46MiJZ5jUInsCArq7JA
mZngLEUeQERY3wSNTP+WWDpzjfYjHc86YTLIFKHroDgitmZO+agZJvMZfA2NEXfK
+JM4DS5YiKxWCvTt2Eaw+f25Lcr5n0KHXZF1Cgd0LC1cbqswlY7qVGu/fXvZYaYd
ibaGwEDoEWfUVKpKapB7ObLNeMJZo1QW+Yis3GfeGGnMqQIY/BebxnMBvWVhk596
EfqWdvlCXh92x/7VUCQ6Bqu3vDIciu9O9EEuPvmezjt10OUV7/HKY7KzgoHj8KFo
0lbExhkbvxX6iNTs6otGv8AHtHaQeaAmFasgVGM+P20lvTXAhzK7Ko4sO4MfCBEp
JNXut68rjuPUFXbqo50th3yyS/Ejh5EYCGelXx7XHmvIQx1lolq+7w5+9eoS4DWX
EfbYUDS2bau1unNxdDd4PDfst9bgxc4oGxkULudEaJqg+gPeocd7vLBfEmYny2fb
szdLzh1aHrRrqPj0UbmZ2KSMs5sPLocLrIBjLUsbwwOTfidduOSaLRAReK7CHpCm
IitlIJymfgGl6YtjZyhBtJ9U95fFYuAhk3xXzaknFhf0IalKrS4FO1mVvl2sH6Md
qQlPHf92709MyFjEUvu09Ylkzo6lxD/r5A/uC1tjck5nigTlXX0QER74abYEgpTG
wFEeR6UL6eEjatUbVPN8GCjHpSpMDCHzicAGyPLkvGQApM8Wv4zzfZ7rjk8PApzj
7PDZuHSXEVCW2FvEwUwIEg==

`pragma protect end_protected
endmodule



module SB_RAM2048x2NRNW (RDATA, RCLKN, RCLKE, RE, RADDR, WCLKN, WCLKE, WE, WADDR, WDATA);
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Lattice Semiconductor Corporation"
`pragma protect author_info="Lattice Semiconductor Corporation"
`pragma protect encrypt_agent="Radiant encrypt_hdl"
`pragma protect encrypt_agent_info="Radiant encrypt_hdl Version 1.0"

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP15_1"
`pragma protect key_method="rsa"
`pragma protect key_block
SsB+fmeIrG2xkVri4/jG1bo/8hwsLfhRrCZLGVt41eM/aL+C3N2yOmoWVOdW91IB
0KZcA2p5VZps1t7NdgXkJLaiInq5XffJKeaMWwPeSDwnxrx9ft94YsTlAf8C3w2X
8n6sxYm8lgp+tPK+mmfv3k5130p6o6GU7hAlgi/hbLLMZ89Q/798FoG+mfrNkpMh
8ULcegUvfS+50Peet7GPfMa1hlAvT/lEGSshbBlRY/qU50+a0W7h66neZZ8cNU9c
7e7tB/zwDA4+Dz9xTItlBBK5nPLByTs5EzXkM3kDOxNobDvYJ5f7YBP0hxvp4qwc
KmihFhtCaImknkd8C1Afaw==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
a6gQnFZwdGUzJxTqT0MpBrvjJ9y3DiAV6eXXRcYuVFsUrjGLTOHPMExa9fj3EWKO
FMv6yo7WD5sGGJSGFg1bVhRDilODhCfSyccugmAgPfV51SXIwB8E4Jparx71+bJA
hfjRoU1QA8AYNuJBZmx7Tlntl7flOlJam0R5nUaE5X/fDfR3jdN7sqTKVvztHahO
oHZ7dJYMN3RjjmJs/TU1B1pwerYe52peXxFrJv5UrI29rqpeVVSkGeh4aJk/IRNh
AM0lqrfYOKYowdq5P91D/iwP5IWk3MCN8su1kQUkWaRHayyWV775g1u8QVybtjHs
RQvbOkjRIlu0TKohJ05XWw==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-2"
`pragma protect key_method="rsa"
`pragma protect key_block
XoGwNgzVz4WiL/cXO6e7jOFvErGXquZZ+1eTtAz8E/lSAUG+ahM4jVXjx98n53PH
p3eVGUraNF/pFwqJjSyIQCwoCAr255Tz1C9M9cOQMuJ6xz7Gp7mcLoprdK35d7+G
7BonzeOqhFipIiPgD6uIbdQ979JofxRkbx3ROIPVPIhnVu5pem4FBDNZwbozC0+O
k5odPX3TlAhI/dfuPxvkLCoBBwcsLi/jCZcXedp04/D0lkI4Ccj2YQ0oaFM+d761
Zk5e5sGcFoubEi987qMaw7A3F0kag8bvU9qwgaZndf/Nu/KmnQ+jNXfyy7Af5i5s
uYq+6WPQEfM4+2CAykHWCg==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=128)
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect key_block
k7eV6obYVAGXNLa8x3++pt943BeRXXARdYg/YO0v0+4Q7/KvugvpWccxknciSTUh
AJxxt7iKNiEBWdOGEk0XCZhE3Pay0y3uN1N+LyHUOgVHMHUCrIR+qJW1ofuELsGg
rB2ONcEifu4xoIAJp7PGMT/reWgZiqDdFbgXgPFOoAk=

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Aldec"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect key_method="rsa"
`pragma protect key_block
z1CKKY+R5LbPUKviofxhUrckKzWDJfig/Bc3p2sM8STnovMFEXEkUIifq2CLohYw
qPEvwAu4/7E/R1AphrvT0zYeMJr8XdTdpNYDqYFjFPZhHqPzOMar4y6GmN+TiYgs
izFfmZ5UN6IyQpsrYXKI8HyYy4oGDCNp86KlRoqbZwuLjjU9W7/7Y8BhD4Wuoupi
cJIWpv5jPdhq2gHGBk2RPE09fiLInoVkUEJ8gStWz0TJa6K2SIu6CF1AFnjrsiec
GPSlB3L6IyO+QMCVlMv77s59nkjLfgJ5bxUmUJmRCul2bQ9u5m2cAprWYT5xMp3e
faQwAsLEmCOaAjwGu545rw==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect key_method="rsa"
`pragma protect key_block
KvGxs+2c4WPwbqaPWy9zAWgiOuN2K+oBNBnuDW16qA5uqB01cztN+MLkKsXVgun3
bqsJe1ytOe5HVEoobdk0O5ObrJZfN60v6/b1uIA8bZuqndShWkfQbtKFbmUgpdG+
fp1ylH//qWLBfkCA9LZHCocE7KQ2mJXYgyznsisliniQFmhsp0HcEA1s+uWpgERi
QAjphITZfHZq9qgd+HT2LMySwgICY4JRmWsGQhwNFBJA42oAGNWztFqSijExyfSm
yy0DfpdPUYDc+ptT5rd9xOPWR/ByMtY50T539k+cSNeapGAqfyXREFPcGMoLhRM7
0RmV/wfIy7hpsd11Dl8aTA==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Lattice Semiconductor"
`pragma protect key_keyname="LSCC_RADIANT_1"
`pragma protect key_method="rsa"
`pragma protect key_block
vumCYngZKbdcn+jtsHzrhRXukdhRAtfEZ5yR8Ex7KghgmMpnBE/wO/Mm6C8pSDFx
ux14ttq0DqCgV3Eo1iw2eKK6nEZS/CAu+qwxApg9lx+Vka02ahP0b92grnjUyaVa
/PBUXimY8Ynam542Lsl9sr2wP56aVHi4IH9DCxDdfmww7vnuYO05/j2Wg5pQ6gBX
Dyt3bNKaOa4LOPysd9cYqGp/emy91y2Tdg16vRUH5ELuRkkVW2mYuXdSITDqNO/v
FyutWaVzYIp0YL7xIvpKtILlYW/gP1bU/GLkiguTWssdcTRfv3jb9QiouWe1kSCI
BgyPjWREnkVh2j26o03M9g==

`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype="base64", line_length=64, bytes=3936)
`pragma protect data_block
NLRZYLWRhY3m17SCN0G7EyyaPMEeggZLCQbfZVyHhwidESuBqFZGdIBQE0a4Q6Y+
E4C6IYMYU+PIfRU8D6DRqHNR57nktkzHKZFJKXrEUrO1qd42uU0IZ+rIGlzmEsk9
ApIlAVgP9STA2y5dfZP6EVxi6/M3SDoH50wP52rQQQu1YfzsKYPzuErvdjP0pPeM
ilo6RF4kQdh+Xv/7VGsHQrzgp+nuP7Rq/RnU++OjVr8ayNhddkSZjeU0KsO1vqj3
LQN+yBIaGPiWfB0gp62ma400mRM9/168+2mBZAS2fq9a7Tz4c7hDNR9cYGfBF5fV
SLh/C5cB7E1xtrwEwbLsMkmMZ3jpH0p/ZiYLy11jxxMtPXy340nxmNLcyvSbIVhM
7A9IZlaM6Ce1n+xoQKZvo6aPNgAsHHOSOhyQW8D4gVpEj5lnWIrfq8k5M8yfxJII
q/p2OTIO20fxXqyH1TRulC1KPPEkZ9X5GMhSLGrMSbyjVTkGzpGRrspdzr3zOzP7
taMITBa9RSOt1CNTx2kG9bOEAfgjZI9ZLvRopsn51/oeuNgg7EM+ABIkx8hXle4a
VfoxvfQURBfKrxOK8gPKjamvvw5skA9Mifr4CvDJ9zURimM+s4bgVqlx2vx19CW6
GHRiNGbc/StxGsY8SNUDe36koQsBLSDoNk2Uriavxsek/FpUAu0NzuTR1Y8W5efU
BQEdUOMNJljYHaADHy1Br9urBnSV9/9CQsqpPOMpglNN2vw3MkrNwsfPEohARLn5
Lv+uvMC+tNK9pLZS2r73p22sYDh8jrmQWf7fsENBP9Ep1k3MOqjnFDtNPDfB5X4x
zUL9+ha726ppDheku8SIC40+gQ0VnYJX0qhohEFGs8yHh9a47hP4e1v+1e4fow9m
Qpbjv/Frn6xTyaUkCFAnP7giNJGqqdPEd7AHm2C6hQsZ4JEwzyl6OWDnq97BzaJo
3pmXV9w2hruXF6QzzDTVG7qJ44jP/tfKlTooRZjlL4GSdvgF1r6tlB1fj6faSEn3
nPRVTD0w9gVQQAdREBAQoEsoDieQndKDRZcwipVD+SLF2oIGbEVM3S5c1c5RSWMU
nbGgdra25s2duhW3CK0PVRux50d9S22Yb9SGyIqzzoAlt2754CzjGNeDkoxK7xVS
xN9QauP/FIxPT72ZB6NlavzxC6qeC+eKE7lbzpAnjKAOKR4CTYlvUEUJy4JzmOZe
uez9EMbXhmsEQvVksb4oXuyiC3+O2nJVp864XTsLQQ1JrTjVPuYppHWcnFnnbINB
aeUxw94b8rIZqUK/gFviGpTTkPDBuGawFXGDiRmk5KquWmrYIe00SWDDrXdhadsI
iqsdbB+9WusvG0ETZU17Xz7PQ3beFuCRxFJBMIzpiqVJEcwEw+DaFZFnPPqQ/Asw
71RsRVD/KiR4ZVLeTUhw3AaLuJMU8InaUcBlrzLTaVRSXzakw6YuyFAC7PTee9YJ
D3bupAA1Hqa0pHUHpJbHPTWWK+yEApj/+dmcDWTwe0Xx/3emcd0GyIJzaY9OlU6p
KQjBzARoQYiRDjdR1RFSNdwd1YkF6K4oMifqO1dIO3PEl+lb4N3cJl9bXYzvd1e1
EpH9tLTshQFyoYOIgSiC5C4AxjAxB5lHCy8pUP6Ix0IdhiLW9WTTvVoIT1Sv5/lv
IxeW2cFx8iJgsXL7lkyUc8XBh+46R4M/o35qib3n1N6sSmfRjPrCQWbr65INOj8W
o68HBGuc+uAFk+Qn0hmdV7bCnSoKQIZqVNJhkszVDxbQEk79LN0iQoBllcdcMeW9
c6g4vPqvzXkH5V0d+bYFn0mb9BXorSxT9QqWbUE9zFgp3+5hPpLX2DErOo5GHDvx
VRFK+2WR36NlonwJG7A2uB6qxb69i6xs1ga+9ax4FSoCdwE2R98iuK46+bMRoRvi
1AtcbuGpSogXrCDnmYLCWw1Aj6o2Kq0gDx0Z9BLNvNENXlpy2+hsEvByiABJ/YG9
gWAwO1QypBkARIP90dD9ok1JJknzttokVvBWb06TRscAIjWxh9SlLmTQyujwzhwY
7z+gUYJoncQYWo6SL2pGX3oNf0cEQQQxJOcvp+tVHHvjKI8m5gtRXhfjh4CgdLhu
gSi+yubnzAuhNzwIL7KUqMB4pTtlnTRQvURe7CdVMwJiW4DPvkpsA7Z0qbCVk1nP
aaqQAl72cbNbtuTGcjo3AmjLSs3gOe7wSvGzQk4dxuJLmPGdOALqPfIPKGqoKxeV
7FEmmyL6Z1hrFZwlHj3A/QRms6PgMU4bm3hnkhosc2dKzS9ita6Yryxc71PBfvc2
ZXXo4Zfm/exwkz9E9tkOkdwB68gzjt47z8FzSoUm3gVKZZ4DB15NhAgYS8oSQaxl
xL14dBUV4+Zq+D7cr5TFj+RsYGCppheuxcQZX4PcSs9XJ4/sao/HsRQH9JAvVtJj
i/2vKsNtFPx0LOlbPVzuPbGwoXPYojHw3T8jrM/Dzc1Jd4ZnLn2enGVNbCJaupez
Kkmw/1w0kT5qaP3jTiKeMq3trBFCvoJWzD8e+0kcBptRmCv8jjoBno+Yfe5+z+oL
L3jX2pev8FucbOL9BU5ssWkRpKx2EfpIGnZV92oW4PfBSdpxcfg6/vXE5p1NVVPJ
8ZTM8uiiY83ysZeqOTsRKzp4RiA9j8XZbWhZFpl1rk/GW7byjkrSEMP9X7hvI5gs
Szoakp3GixTwyk+1uZ+FFg/aw8aE2OuDm5nciGxMGTQm8OyHVhlhbAPSkpZGUXse
SOBHv4Ara/Z86qhNuSgYZgr5upNV97cmg+UfA3Zg0IomAUPjT4Tzihtpcx0t3kIE
shv0XDu+JeO1k8k6zNdlOkP49IrqX77ytPNV9t3y0JXI4I5VJX7fW0bNG++uOTOS
cOfHK6LDBT7FvteBf2/4aNLDnDtUZROq9jC8BC8IXwUKVUAArLkU/+hojEMjryZF
vKrNtXPLBlQw4rU7xpYYGPMD6RJEltHSHs9NnyBYVCPd5UeYBN562naVR8UgY+5H
z1ybOppZryFH84Mt4AGCVjzT77v151T6mLYXryUXxdfsB493grMpQMcQppOuscqy
6B9O0UhYxK+ySX8qLWCL/8xtCacRhOXpuaVmmnP0TEhBVpRSf/sQv/nkUVpBFDz0
DVuBxswijU28GjIMhVk26/+Mh3N55bMjzAHFdf7IwLVCLxbe5HYX06G8qH9I07uM
XQJl3GefpTgkWO5qmyJ6zENtK1BLmJ6Hr8s5IQV0EzImHxsoSJrUdKFewA6xOvpm
PaKTY0UYhUfqGVdccvgSwjFKhlss8WtPyiCztxeTP0DFpQoYVzHq30A0Jz5QMTHN
ADW8QAVOfNhsWSLggLm8/z32I3B7VI7fHFKYI9Ir+getP9gVKKG63lFAqtWdGqMF
tUzaTJweR8IDjKE/yImUpDRZf1Vh8WzlLMFMEHpVU2kGurEmEAOZL3iC5GcJKtIK
or75NmBw0tA5GCegCOtSGTHAY4WKbqc49TJchXu5uMTCebDNmMVwVWqT8rmz4TmR
StZ/Ya0+2wbGMY3n78J49f8eloR7uLBbRrxJPgCuqMffq3kYwE2woz8OZdMDwBen
UjmLM0XXghqBtWC0xT+xdPLB/jWE27YNKxnHzwCUYTOjjMy6SWEwi2FNLsaheXRO
xhBtv3S4gIETXZEy+NiSu9mxhKhGePbh94XJhEEVC4Pv3934tYVyifumZEbixVK4
wghxmg6U7UbpUS6QJvXR2ypGqwWBY1CAlS7rjwLzgr+yLiCxofhE9dgybpinD5h1
uvMO69ftGH+qTWpXbsa28KcehBeRTGBDbrCqEbA5WrLyoyYi9nPpZhLNoxbP0IJZ
5MKCqTru9/aPRfeQUAKg6womb2lSsnyTukZYoGHXjO9cx/HeFl9eTk9ENfdE81Ox
LoEAG7k5vQWyKGEeCEJu+CpC/3/w6CjK/7sKoQVfl1f09IhA13x/OLNzjF2QuGzE
2SBACZTbo+kBvhYgTSCSR002/iGeoWyxl3utuLDrrhg6TCh0OCjncI0Fdqs3AlqG
+o0GswbxWQ3QRu28L3WPFG8TrC3+fxilI8pN4fsHNJ7K1Gsf/hopcmP9zqYUuiw+
IMAVmzh8iTg4h5Ar+65aMd9JRUikQ/oCgJxGJqBHdvCw6B9V6D3PIyIIK/BsUiVo
dbfhUCIkPH9MbQluDbC0C9FwHnCJLJ9UzZL/zX9QECHbSae6R67ccDjW6APFHY23
+vGC0IGN3N4pt3dQZQZ+9ssNQETNmRn4vcUjBBnyYVjcpEzsbvMFl66RoaYVXnuz
rMMZuoLLcSkt/YJJnxf/Z9EzV7kG6qTLO9ch+NgHEJ9PBSwHIRzkvA5j+iXA2Gnb
q6aNkzDlu38cuA2BEaBPlmYx1SXXkNudU7tOMFzCQCqJ7kC6u9YvpY7AwDSjMcWL
kHTzCleD4LkTIrdJFeSibkuqDLfFmTwEKqKackwBjlWMoyz4Ia+e3+N9iENBXl+T
S4wLMy535upnJwPvF+nWepX1tjV3/ike2zP6/wXBuE1TVTfvbAlpOCoh7w8PqJpn
K2x1rpF7YYTrRjm7X7aDzYgdt7Ya082/mQkrEdypXffi4zrcLRoPd0f0ZDzESfcY
vr1yXWQKQKyhCAxOJZ5/Gq7DdnjLXetK2vFf9GL2iwLOC3/5BVKRs2sULiQX5rkF
cwJlymq8LY4W9xsVhxnKvLi4Yo8ew6WV07ZIXAPWqbMSvX9iILevoFt7HaAXkW5l
2qZImRMEvk/LULPmNEMHYUFle7iaLC3SBNjsuYWAvHEgXXrOtWafXsNa3WbIhOQ5
2NT+2M5niaTUyQLXlJ5Mqjh8ySIK29d8eDNp5vc+NredP1X8+v5RW3NuDKLQrSIl
m5kwA7e7mVypbDss9TmUP+3Ooa3oNwXZjUzog+bz72HN+PYVEK1hUnGuLRDJCCek
dYQjbg5EovFdfqYdO6P7QinFaxPr493K4V7JFlq+lA8ENt5QEWDrMiT8ETrwJZPO
lYPI5onal9iqIV/2jV+rwXT/acaksWT451GhNVH+6FcqtnE2p7H/QYYiBroFkgMB
lG/X19HO7pT47mpJr8esA4xNZlX7TtKCl4gTpgBv7ANUY/hSk8jPmAstaz3Ag775
tAQPlrbBVbElmaKac1AEM78BoDxka7+7+D8xddnP2aAAyqEMtQpgN9/rcJwSt719
I/invTed9c1VzV/GXs0JWvSiILhiBme/rZF9oixIRd7foMz8Q3z676yzrsclZ3tG

`pragma protect end_protected
endmodule



module SB_RAM2048x2NR (RDATA, RCLKN, RCLKE, RE, RADDR, WCLK, WCLKE, WE, WADDR, WDATA);
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Lattice Semiconductor Corporation"
`pragma protect author_info="Lattice Semiconductor Corporation"
`pragma protect encrypt_agent="Radiant encrypt_hdl"
`pragma protect encrypt_agent_info="Radiant encrypt_hdl Version 1.0"

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP15_1"
`pragma protect key_method="rsa"
`pragma protect key_block
iM05l4Rop2LyfJKSO9xijou31UjGwEoIVjrvtAx2QZFXmXL7F73fabugaFVoYGnp
elkE9QYCO3dO4ncdQ5knVxgfiSz2iDi5fxsRV+Tu8JmkPehw+ivFlCFGtnsd8iTW
xrKlmilDr1ehOCx/TfSj3lX2Oq2krpAiuX96rTCdkpLa9KlKfPCDzJyJrx00qcyc
PMVrnSazIhETVP3MUYH138IHByi9RL2fAkL3/dgNjHA3taq9AAgD6bn8JE945tQh
vSuCxDSD6N9IMsgOgHjcXe9tUk7ZttwZRfO0aPlsZgwpLkLr5tPm6ZBbEtRgNtCC
X+kAQwaLKUR6jffu4XVIDA==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
GZEr5Afxi36zH/YbXldfKTFVXj9ea7AGGou1F1UWPM600rTxVJgmET7CmqfTxMIJ
wIS0C9QVkBvtqzpJyWEmT6fAj8rH7Y3fuhYJ/klxaRMW1tMm5hgP3N04+C/1JkFT
adiyNlHv2yxkYiZlNSFCZYCHW+Jrt21hNrtKrXxuQZmKoAazPoFaBirtqzbz2E4C
S3dC8BhJCDZYY2GVFTsWAciEM63HwcyrdHW0H5LOpqGAF9RcDsw4ACFESNJdqdJv
2Kl0Vhk9otmRv4bVCdI1KLrSzDJvYGo+EvbnKbRT8iMkV8oUH0AgIkBcko//Mfnn
vRa04/Swg6hObOPGgXvfNA==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-2"
`pragma protect key_method="rsa"
`pragma protect key_block
oEfM8HEGYqHgXkv0dtGjfG9PMQI5/XkH0iwHE/HR8r6JijLaEHEhsIen2wvQHsNx
s5IaloBrjDuTgc2t3C5EGVWvFBsqZ8TO43PuYekjWcssyf2f+ksOKsgYaM4lLtso
25LIIDfWlTfj097jvczxYtR36xl2SX+G5BqmT0lYNpUG/OH5Y6FgqQgZa23eM/iD
3M+TvBTlbAzaMrRzEJfejI7dv/Bs3kBQzNGVUx20ehpLVC/z3LSVAhfcJ53qXjWT
d5H+0ov+JTwquVBMB4CQrD16/bcDLvxZjjah1yJReL3BDv5qoTEwEUoRr6XfnWnr
febsWfCDCC0DvugA5Xqabg==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=128)
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect key_block
ssvvSH0f253SJvt1IbEOkWSB9peYuVQpXPcqYxQ6IgzluNiKGGBpfrVGqqyXtoHp
ljysFm6nwGiEzUAub/MkZzqMmN4XlL34wmG8JUtcWB2DY29YeETPJ+4xemINEY7T
sc41xzXdaxYagY2B0SLXJMBYgrOBvvQjjgh3sswiOy0=

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Aldec"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect key_method="rsa"
`pragma protect key_block
L24Kg+zQCsIlTzcYtm3bjq4XLL/PqP8X9Urf/g1u/Coy8yhA35GGtPWAWXX3h79y
cQGuhA6q3rJwQtaNqUoBXjwgGPfCpEItaJvoH9UMgmvyDOSnhkLO8GfoZ2YBOTHP
7ZLkMZ5W7fIGTc0/HAMnM80fvcmPV263+9S8+pjbxLfhRFX8sTZ/cfTp7VlYsmdd
ER8O1tNBO0fAT1FxsehRDrXj7tV7/JFeM4XIdJadhwK40vbAxp5ab5twsSvw1HTx
BjBUT8A70g/JdiLbsqIgFJhM42Bmvwq8dUnePUdjXn6MRv3gkxcrwIvptOmh50YP
CHX11ikKh2bk47jkeWtzuw==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect key_method="rsa"
`pragma protect key_block
i79D4qdPef4IGwJw/u+1bpyXkGvzf1aTZVMkmWYQQmqHaX8lxz0mG0AxJ76ALzn5
fK7cTQ+mu7v6OE5fv9FG0pfx11WkCuExRVkL3T1M9ysKEuXYLKvY8x2IDREXRmzy
mOU+viYoSJXI10jbptKiqlNzBlKIrBY9a7Suly8kIB4n/p9DkLx8TtkMJcqPW1nK
SkQWb3e/9IVdgqB9YN5V8qUATib/FoeiJg4TpxNjqEFjSFUerh6Ddj2F9Xipc08A
IXcB4rQuhgGCIbDWDVY4A+d4V55Ga3iCD/dWezGgGM3TqBRmaKXPW75a1JROmDr6
qellOYozRK5fHYeNM/wlfw==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Lattice Semiconductor"
`pragma protect key_keyname="LSCC_RADIANT_1"
`pragma protect key_method="rsa"
`pragma protect key_block
hx4PXT/enRolIRaOchDmZP9GJPgPpU9Dv/vosHn8SJ+A2EZns71+rpdZyuqJcFjL
k/33W7hJvxuaZ3w0pohvppkWNrQbmE/GCTe0ww3C3hDRAFqKYFeFk5ZxdTBpRdvF
vb5lxn4B4DwXbXagT275yjt9+VaZsIuGthCRYEv1v72sanWDpz85fUHrkfLYMCRv
LBJ4DWpLDHWiQc0KtSysYdtNQBlpf+IaThmshTu7e7aeAjmgROB6szDbLFEAvU3y
qulGj/nTyD+qgsDEXhFdaEqY2Vychwh4sBbHc02C8asuFNyQTuWqswANF0JpIWqh
RlFZsgquTGQCplR8Zia7Hg==

`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype="base64", line_length=64, bytes=3888)
`pragma protect data_block
ZLo6XclzWLlqK68+QlZVkAxXH2S9r2ZEdJ9zjoFHTR+WjSEQnDKkgCZK0elUGaLy
zYwXvzg7UqYHVrJ7Km4HkrcjOd6peCiyjcnNBGqMa5DL4gJNpp/32iZMdAS/wxfX
P7YI2DOTWJ6BSZNibzu1srPGdXzVnB4h1+c3CSS+eWO6TAPMoWqDMkd2lCFtZUz3
oQCtGD5CvJeRXGjRouaMjXIrX3mvBaFzQKidt5Ec3CCVFOB+a83KohDb45EcA1A4
dw2/I4NFmpfdtLApw43vmwlXS1SpZjyTZsb+xFECVf+VoHH5M3vH7oUVl8x48Rp9
P+4KQlPo/0Bfm8/DMgJO5wTwZDVg4/sVD8LxX4YoLtLp1w0y3U0UNW5V3XFlLyS8
jhuJGe0cj7+uDN1BPc2DvWlLKXZasCxVewvPUMchH0Se6neAE57Zm84xY7SCk59n
nlH3nukz89fZgg+v3Hp+QCX7HF5cxun1QVkw6JdoTEYVwLu5V7Iy8r+D87CEZ7X/
PAbI7KEDbsgpsuqypQftDGTjc5bhbDfXyN+pPVkvVkH9ynoE5n7aERUp2a/mNWHB
X5lXGZKpvo5XedFeW9bK1JiXl8yF3ayOB9dGlyTy4P4ED+KLNPfkr8wKLmXSXC7o
v/7LqySwbmUZKcjWcg91mlUBmDRepUFofm2cTCjT5lSNdBWVeRhqA9r86QerF3lW
cfApaEOuRF+zoCK6xtA9vzCgZAUt4Ia+2ODom6KWB1/vpJc7WD+CgUdo2vwqfaqi
2H3MKgQIvBMnpCiZDLVs7Etj+ObFqQznIl5Q+1Az7J4OWvhMfhLT3VbmIQtE7WPL
F99lrWMN2BprNw8EqHRtYuh+gm56VT8fHaQ+epUNyG7Rt4VS4q1tzjAZuuKAi6cS
Ta45vmf702cqXJaudglobmeMWu2D3fAuLQWDa+0ucKtGu4uHWgMCQS4GJeYqqgHl
5T7wS//0Rpy1BINfvvOA3wym7yO4fo/PyPWCVJHoU1wmpncz/C6Ez4vPVLP/NIMR
TPcuJfH9v2mCU8pSAPYARbZaZv2MXE1X4+Te1AQoM83jJ6XMIN8yDzuDArnpLqcW
eck2vGTh0VXGe0bB0OP4SPwoPHVdcu62r3Uq3/cQWtMVUR3rwpzyjHNbzPNLqNCX
XciY8FI3kFiIuyZr8wZwpHEMb1DZSu+4wAc4UdksgSzln8w0GSlWg4KC80+/LGtK
oLsB3GELZtfKw70N0G4DUeBDDmf53jsWNR7Sbmb3eq1U7ku8h0HN1bIxoz7a6MVH
sYj9oSOJSf+Y5uAxQQWJ1qG8oUo+wJEESFRUNHFV0uSjVnv4epGzkZ32sNdEbtOH
CwO3WtLt3/t3cLvRbG/FxI9W5iogsormCfP5VtVzaomy0QcVqxFN/H0Z95rGZxUI
Qp1AKNJ8frYQQBo8ageSbB2iKTFOI9fR8jmIQ8KGnWbro9M3Mktmc9YVWXMt2XGS
fQWhUC3y12FDHB3r6rk190+uhaJmOr5LknaIoijaz8s9dPKoC+SxSXQByymw22nH
/CxChjulAbaxBo3yzDC0WOtQiz/aAPRa1uPVHb6MS0OoPSXE/P0s3bxaxSgX5tTP
FuGEIhHuml8wRPipzRncKqLGkcY7UXxXjfuP35p7l/efEJBTTwokZ5k8cTUQBFTG
CeAokt/qnhQMV8KXS/U5zDLAG7kuxyPceHtf0yC6/9GaqZqOnpLLMf6wEw5TB2/b
bB6/DdVrC+R5i8dvl+MzvK48Ij+KsDxKTJ7igFIEsVH9EfWNmG4BuHQeWpC2JR3Z
EFFNYBsDdc35OqugYLMCg9sFoHra1M2uMQhs64cYBcKfh5ZOck6Q9In4oQqQrtvi
n2MFj2xHeq4wCXlOGIj11dtfeG5FFoFM9m0yYi9N4/RjMJ4/JZxhXBE9tltyDgRZ
2fc1vUya3ok5LSNbok3qLFZDY+R7KvG6GvvDBjO5wJmjMH+kGdlRlNHzHvCKJgiO
FF/JdbgpdGviVWGKwY7L/4B9qFxeFIZQ/grIilLp8qW8lxdqlu+ZvF9amZW7Sb6V
7RsFCT7OSREho0m0gmDAPNV+23rP4X6dnAvJ1BI+X7iHj1BFKogFTmAq4jQhXlwP
YfCdMW6SdG6CGhvnCA0jYpCfdmyBD4e4kc2P9+UWrRKF81QrzF3i+8IZvW/HA2us
tSR55MqQ5TUy+Cw2Y5U4YsMIb4YLfOQMBO26zxUONeeFBLrtIYwGB5GeteaFvLQ6
k0Hv7pYII4lme9vN51OsLbfGTv79bSyMhnDy3qRG5XxSqx32iSiYbbUwKQv6hQ+z
J9FuWbBnXq0lhiTu799wo/MhQ+5YMWzr9QAOdEcRaj3QM0OdF6Xy9M9P1W0ZQqz2
585oj0dCru3Ao0zBhmRDYgeKV1clr9ilw4HtXT3ONrf9gllW7Uq1eh6+8MtkizwL
EXmMzpk/gpmMettBbvCzQX57w+7A8GJILVvHYFt+xAaXg8kln71lu3+7oC9nN0us
AX6AsQZ2YbcnVJ6QNJLPk6ZQ6rqgUxDh1/hS5N2KXn+5uhHAjJOsx1Wo/ODxqF9x
6aPTjKblG586aU4e0qHmWRIYNvBExOf6bAi2ctJY1MBZEIRbkHWNZNJN2f5J1Yp4
TlrYTG+Gg/QHNlKtSt3IFN/N1QIpijDD6IQPQr4AbbJgLzRFdCYWIWwpYtO97Jzf
u9mbcQMILsXb7n4dVL6HbW/W4Cuc/nv6DDx49harFVnkyDBakNsiaAA4y2mSUj5z
sZagNvrsrp5Tp+eEGsAarjOmENP+HiyUF0GsAzdNAKvD5ujdtoOA9U/DZzTtaw3S
TY19yy4mwbkoCqsKzEZ9/XZdULZwWVYAjvwK1QuudUxOpM+q98m88yHYLNMvOBr+
osDzQ9FNrr5I7z/uO2DpzjffE3+k0wYNcuKhHLD8ZhiIhexAN5dM//FWdvvc5kI5
Xwa8HmCjOwhU9A4Ks3CsPLSPYZnS0DHb+ckbBWcUxB46VnYdX6rzlKVmyjTr+sY4
xPbafvHMt3x4CFitw+DwhN2sUgPW+pnJtHo5W28H/F9Y9HXQoaj8v265OzmEfZxR
LQiBppnjDoUVPN69T27y7vZ4fqyD7h12lOSJIVVExAXm5O4Hkcw+/U6IpZYNCynz
90u4xLxYJOq7qlDN9x+bJB5HqUXF1aJowd+dssR0Nun+2eWyQvRFNlkdvQpz9I18
pQcBD4kadeYqS7ARexNU3HGfzjPnJHZC2OmUwXLXhcfyne5QSv7OFikiEQgp8dtA
vPMXZnL2Aca6SWjtXemG8s9Ll19bui6xJW17bN7x1Jsg6UWS8AV7nKMEx47jWO0Q
HQ4opHxR6czZQchq2/ZSIEVOK+THLfjlzpMbHVmM4GsNWETrSWIkmJ2KBLCKlf2v
UIzlr0fHNX97vCHo5EltshT8we60E6V/qcvkzJCyAeazcYFWAhG/Ae8IxpcjRyqC
7/JPYp3lK68hQ8wHyQJpvjzErrnrvmwd6Y9zoo5HNFNMflHMwgYRp1pqp047plRe
jrObGE44yDF5ZoTC9qa1HItUAkvW+sFxQq6s+q04uTvONsr7j8RFV/+UpT3UeK+9
Z/Lm++YTT+toKOTs9soahmjhQPSbfiWJAeAoj7eqkANgLPtXpNdqvfyY5O+nAaB+
c+EFybivWg1/Tnz3mIQ7p7zWd2Ldj7ztv/hH6COECCwi5c0WknTqKLKWiSGiufDz
OtDgpPnqSwgGv5Nk71CEKVDzhjdidDBwIDntww3WjmC0PgS8SlG8DUlO7hKLAnkI
zPZChjCvdUMIjS35y4czwM2495mQT0hz9jc6NT5PBXwp38UKtKCIrzOAf/NyZPWr
6MLUxwL3Y4K4W2v2ja6bEx7jPREXHoc044xzd/xPM2/VmTvoZ30Xj72n9G8WHKKE
8u2prYOtm/4uBcnRxHG94BlkXIuPj5nJhppFEgcsr1AXf3bxn/dQqYsorlVAmtk9
wAlJRePmG9J31kfi84nRm5uuwPNSKUDEGjxV28enz0piQw/in6DkIGiz7eRZnRiq
4j2+OPN/YQr1htc9JHAaJyI31nIpwPGwdIovDBCL90qZkh0EGoAQpd9ECfPTlEed
AaO/7Curgw0+dAPkX8Qoxfip8wLEXflGVXtcec091uLNZ9ag9i+p7gEv2tymRbES
nOoF+iZtZkQ8lqzQxNMPO/jSSJnvt4/xIeS4tMrspTBGDcltEjBeOdSYbxBpY5t/
S6CcgI15nmHMteR/CyjvSp1qL9eTNl7O5wynAw4Y3Ixh6GxRY3AG2U1GTdXL/upd
yx8vLyZt8ON0RUlH9ed5WxtjtskurRZSJTPGlkxJ/DIFxohgeN5fGmocpiwD9ZYV
95tRwQ/bstkhCPU2+EH+PJQ9N2cMOCDdY3j5U65NBUT+FgCLBvrdrE8mPr2RMfQ+
0+VINiNTgCOwnPWgm5h8BIjACyYrTGWgKLpQPtljgLOTnZpWjepbWXDwA55sHLI8
L9r+StMuQG/yVhGOjg0wJzhGjJv0u+KCoI8yzWX3hXqTGZccqjUmoXeKcu6aJ7E/
Y9/1eGO1KVD6SSlIS1i07BZv1HCgXRHgsdmCxJ2AUUwYtrCB6j2Aq0L8NSIVc0fm
3gOFUhkVeTD65TA7m9a6QZHIa9rAIdkkHZ5583efUT8bN2Gdd//Bb/+ZqvvK7Qot
hkeB8esc66QYd/7QC9tr8jRsWU+G2RmVK/AfQ6+tEMOBm1VwXiwo/0k5aG1wLJGg
OxDbLhrpqC8V8X1pP1ocYYmLvGCT5IntxDvqI2TmiblKPCr3fwZUq6POQzYRBECm
ymEW3q+jqNjmZp38yc5DJuEDSc/i4HAXIb6dy0/1hBFaxoCf7wrqF/Wxa7rXPdFG
fPmd7m9026Lx+reX/R7SRpg/yKb0q+O5vZhofKwwc1aKFYgKtomMhyg6EormhGkO
pU+fPXXGX4qYysSpN5e7UUE3MV0eMDeiFFWG9x8rBEvk/IJdWfY54Pz2NDtaliu7
AqjPXE31kYWuSqV4L8cafoc9XMMcDe6gVnxRsISY/lfo6krycwwk401FY3ylnDuF
8rcZLhgDVcVvzUQ6bKkLcomOCo1Y3IOHufADtrW5ruTtIUu3ovyakbzGrw1lHGdB
YKhNkGW7KgFJfHE+Mmg/qOBzq9GKOFx1fg1e3EtgPFbGeUmlpei/sFXqMM2NaCVW

`pragma protect end_protected
endmodule



module SB_RAM2048x2NW (RDATA, RCLK, RCLKE, RE, RADDR, WCLKN, WCLKE, WE, WADDR, WDATA);
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Lattice Semiconductor Corporation"
`pragma protect author_info="Lattice Semiconductor Corporation"
`pragma protect encrypt_agent="Radiant encrypt_hdl"
`pragma protect encrypt_agent_info="Radiant encrypt_hdl Version 1.0"

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP15_1"
`pragma protect key_method="rsa"
`pragma protect key_block
WygC0ziaS6y8o5KPt/EBBcPpwiK4UtauHgSqDXh15TqEvmV9NkPvFADRGk8RlMVL
yEiP10AGOX43qOIXGiS91YtG//8kHMaG9iQmlshFLG1s65VMp/BIWtHhPxO5DBnn
XIotzc6ssPq5FqSBM3UmYlXgvsfupccOUbsX8S4H7tppT1pAAaBZWMJIFjLuFVny
BZcRkFOl9ShrG6NP+Lo0tj4lprul7UwjLMJJOE0paYMtWbX5c7LQOsQTZsZuml+9
9v+48wVkzvVajeRxtSvY0G0pYGLGRuLmF6YhzWP6dZWKTb/4+wJdl/nJQRoHmG2h
R05slXzXhGkiaHXnEVJZBg==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
wmeFuPjQRVVYlUjvLbiYslFW+GFLS8M8Ac2Rst7KL53a4EQdPahUFNJdDrsVERdM
YshNIyfEFa8GVv7JlFCPErStgQsIDs0bk4RmF/ad8KenQB4o6aOcaVZEIuhe4ksD
veHSe/c6SpF+3oS3COUO69S9mTaY3z6QgsF3fq6WX2wFa+TSxFnPC0v9SIpCmRed
U+wlG0Mm7agMbqm6RB1f1DeUqvPMMEpr+6V39/c3kmkyRTYJ+yxO28e46bxn2A42
s1HGq3HwxGb3NEo8hojL3egWQGs6S2bon3ltYAA4a6kUELSjSINeSk5RX+GWDAor
l6qOqSglMySJio4BkY58+A==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-2"
`pragma protect key_method="rsa"
`pragma protect key_block
BjbiHiX06kQ4Gzi2hX/Eexfazd4KfIZzUsc6QeV6TCI72p8x6qDbDqsJxkHOqzuJ
6FO6owGIQpBp58ikbpG+G5/gaVrCE8uKtw8RR5sqAXI42Y0dsNs1RbAlwfDSAweK
t57o+niIzwciu9pWBvnsC4S2lMbIoqFimf5vwCfiAy2jVfmhS4yd3GTq+ZMo+CEi
2add3POmOp8zcTxaf5pXPVNkxxFFMEoH6fz/4MfbpVGwB2MbQbWY9q0VxnjHU7gQ
dpopkAvCGkQKjfUL1RZXrDhIJV70TgO4Pdu1yV98xxqKayYN9CBGbkMk/PcHc4a8
rHFzECjIx3yrFLQaa3gJeg==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=128)
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect key_block
QSy2QQ//8oe3bP2QN2QUDZxgprdoLBaVNUh5tGPrNpAx20nHhwoc8WACFa7715xs
PCDV9uMip5R2mvEi9tK16kuxklOqq7YYyXskZVNO/hHtbZZ+Va4MfcXEEMX9M1qz
P8cqlUQ4xWwXWFyq9oEpMgfjp7KprH3EDeAiyXA56Qg=

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Aldec"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect key_method="rsa"
`pragma protect key_block
KCJQbDzVo84wHAluGJcpvsGGyT4kSqCyb59NZgD69f3hfb4Pp3MS571/qRU4Wo8L
YDwsCx4qXjr3clQdUDhpoZkZXYa+Mb1qclGhTVaCSC4vsEWSXoEFwtx0PIzyM8BD
KwbgZGz0gmSEloPny7RuamN9cQ5XUuS1lsabtIp3bYbFxxd9N+GW2b1uhtbtIgpU
cWA5XAJG9VA/nO04T5E1sjszQPl6vuQN16J+D5dVGWFhWAo7p+xSI9uQRdYP1sh1
2pMWnqlLsfLWQdbvk6Im/Le2nI+pCR7t0FUv3C7fDJr7AF64KavsivD4Gb9Vow6o
cZ9Xg5DqTCYYXytAz+VUQw==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect key_method="rsa"
`pragma protect key_block
bQ/0MwfsabqxwDOawfQRKun6y72N6lWl80n+yKWp/iXFXCxvYEXUzp3F0fLs2C3O
2F893bnDW7vkE4ZwACLJ0krOuXtm+HpkmF1WXKgEaY5xaIMUGWWMlMvN/91Mixi1
JSFVYkHbTi5+kFGYLUdWWW4smP68kkNygUVzi6RJZ66beoLV/p/tX5SkXtlic8qO
o44ddp+nfHQ4pqirfIl4lm4+0ZBeYvp9g6Yc+j+NchSf3XQGMp2GlbjHGXWSWdfb
wY8/KtxnLKGJDWTVM81dZMsNhb7XzilGcRR+VnY6xEy4MRXceuNmqoq5roimnTH7
+Dyhez9mWvfOHHPWx+kHZA==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Lattice Semiconductor"
`pragma protect key_keyname="LSCC_RADIANT_1"
`pragma protect key_method="rsa"
`pragma protect key_block
Hb9tUwbwr4Ezv56IFWFSVXoRaknatl/sz2iDU3xF2XtgwYPjmzvpf7LO3i6wVUHU
z8jpM34F4w1JfjsRJeHF7OcM71vnZ9F104JLw0ve9rqcn1vnERZ3LMmi8JDTTQEr
08Jay2NIrua6jAXtABFSKt6NHWFBBPjP0WMMDvmmlL0oqR66Bxth4M/EiADfjMrd
CK3wU6NPrmyFPbc0NfGsBS/8jylW4OS3kAI6hHlzK4bpthLnNMDIb2zRWGN67Ik0
EVzPpaNc0z2jPadDHS3ExhMWAIAWopuYNADEEcluzVMwoyUUbJFeHkX9s0JlcGYT
eoGEzXh3G48oeh/t5f03uA==

`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype="base64", line_length=64, bytes=3888)
`pragma protect data_block
85mbbTuOP8JQHhZCS/XLBN4gvsS0vcAnCWkTqZunAM0cFzOCV9yWCspZAIoqoyrQ
vJRJBBPzjtyEXH7mBB6gEVJAUf92WpBB/Dp6yqmDUrp8D2Ke+dN2ANXWMVj0JRy1
6Na3TCP46Ly4dU83W7Vk6H9za3PiWHcpBT/JMzNU41MbqUKMNJRpb+c6wd1j/3/x
6p2px4jtGWafeS/xGoQ0ZJtbGrl0Z4Fl2VpjZWrnEIR1wGlRDIn+6jKgodYqoaf8
EsfhBJC9okZZ+zhEzKLVvjwRvC19yBhqXoKJB5Yz2B8jYxZsVRDpOvwRHUKstY0M
BV5Tqn5HmZes9shd+75EG0WAX1X/6pepOu5+cyUtVT/xkr3EKp+0NMwJHLkmRH0H
nBW5xQtRHZDS2oyf1oFq4tAnM6Yc48jvjtnoLeTcr7JB9ytr66NdRqcu10tf9PwJ
q8+NL6sAb2ZsWHMN8TpyhsuLr3fX6AMyYw7xGgoKEdGu/6AUAxRDIVWaHhz24LhI
3t5fzZsQ7bd9meQS+kACPSHq/ehiXw+pV2GR6lVZFowfr8lYwRJuqE31IZAmqfBh
9NguXnqQtBY3/kF7TlBxQdcEKEMz7KBqTOXWmttnZUTlGLrZTJUn3+Ha1C9oa9Go
jZM9Y2Ita+QkyV9SWVQkJUZAcu5fIAoqGPxkJXAtXqfwMz5XTCODKoNmVWK/9vob
NfvEAhZGPDDegD9xonsPSZIGNuovHi1EpGH/bA8cbPhLi5IKOjw9C6Q9WefCK09Z
VV2Cj4xC4D47np/7XkDjhP4jdzA4SDseErIrMzCFZRQxmHby1DdqWZ5ePpqohWtK
Agbx7SVerYqUu+csoiFfUIa8LLr7PIGj2GPh1pa2/sNTW7+FSbR5bbKk8BAwGM6H
1wSZuLm5GCVZWIx0z9yXZxEI2mnySDV1V7jPoO7HhcSmoinJjURghqX6YxseenGE
uABo5Xtbt4LB5KQ7QcjcKfng511vbB2Rmmv+1cHl1wSFoTB5abcXbvwPPos8O4HT
dH8Nb6P/uRx0iILMMX5KdJzFM+ejS+ZW4NOT0ZqJXVoYLmF9+bKjeD5vKTQZEho4
1jv6IsZYMBf3VPsums1Wnj5RmvFIWRhldAydHxf/pjlma1FgbSwLezvViMo/50Hj
MP2hZ2SHUCS9jknp/5OoVYLklwqdrQVHM22aZ/m7aDzsczYjmwW0PPsdDA4N20ep
F4dDKsu3ONMPXJzof4qD6DYpe7Uv99RQIZ0beeCA9f0c1VnZ1kyC/GDMdUK77U75
TyA+4s+hJcI8xTvmbpZHyeYOV8zT6DLTGP5tkUhO2VHE8OnWMjIUD7pf3CAmKXGO
m/Y5NssluWpjc9M8X0tl3Q2e8pljsV82Q6YUstzw/oTpMQdGNV2b/uuA+qrUIy/D
Z4w2S7Hc9lZl3XHnHfK+FJER3Xm7kFSfV6PpyUmKl7Xp2Yw7TLAtiROJLr5gkW8B
h2ALf2Ui+NDEzJyFaJxKDwMMdFwYqDWnJoLuGTTX+3VIf47ydFnnL6rofhK4WPaC
1a/oS3tYdzCnsm4+YflaR1MCXdMJcEkmRGRgZK1yjgyBYxGDxba1Thv4IMrVim2l
KMGg0B05vOC6KofhtVyiqIS8DuCSSH+2VfHzJkLUI70ompmXSGpzvAfCCW1aoNZz
vFEUxELUMvFfk2lYEtYr9ojGNVdY+09+KfY1A5gItKEC6MCbVIh9Mr+HJNumLR3u
5oWw72gXGblz7w6G2lZIlmfYZKGs9KLd1+98MZh2rMZzANoXeNQCgy0BnWXeMLFC
314Z+wAehAlxxuzO9MbaU6ctDdDqTlJ+NS+xeSeIaKXaEqRiZlDnV7Rt3ONtADrd
EMKdKqo6+sVXINf9UNjjZ99lMyE9rMTlE9/+8Vqnn9z02ccCTOgWDAQXzUwuAltB
EazpJJEU9f+PThB/sIiB30+TmoF8BZK5x2JbdrPcMovouOXSmmD3cr3ZbaX91dXZ
m1eZRXa7gC8ReMM6vkPm2TfwQqeorFrsUca/gmq4yV2Brg1e1Kr2iBglIOVYYsRT
+EKW0kc4k55itdMtOK35VwEp92EHXw9kZguKTZvewV1P7wEx5Kw8LcEQ0Aohb3Fx
pLGAY7v8BJiexY6x6loKXMD5+7/Ms/BX3TWDfyU6rLH5pdxmHfYisn9Oyd2scG5y
KZZ6M6dYvSKnqvx0DsLi8qZlIjTQFyL+XspJokJ2W0bNfyOOBsXccn/XQY84j7mg
YJRa16VJuVikaQSUuUBZuB/tkQziGRDhUB2DY2f/9DKVie5bxE5T4rbfSvhpd3+r
Pq8iUgF1mEITiYiIr+EBCTcACy6kCsVTLyFh97Ef3xY5ocl49Cv3MW7suwfT8USI
My+0RjHpT0zxutgYj9mIf+4/jFIkS03wR1uwaEkjkBECAztMgO0qxtW8sUmrENsV
BLhVmK5jNBD6+1YpiE+4UXlBWq2hF72FdQBParIZtBl22AHBryqGFKCBVH+p+Z2O
saf7BLZwEWWSYadRrpMJ57ISFCfZsIWPwT9NmmOnpRI39jZ7uB0DLurV88fQtpWe
zduFF6QlJxvOnKjGYUobxe/OGVzeHaQSLO+HABErngQKGOPKZZZ2/TZhStEnJ+qB
12jaMkdhnf890L4NMwoCeM1dRi6R6HhgAvwvJqh6yYoASSmBck/c82Nkn1CCuA+Q
fZOp5/UZkvEAtOY3xsDS2mMxEAhewSib8u4MedWH6Bytmwy9q19jXMlLxDb3FZj+
eyUFdzhrzPAk7Bq5E5WumX2E7y5ErQO6Z+lic5VaFomnabmnuRvC5dyBpMGgVn8X
n5RxeIeclzZeST5mOTuK8k+NDQwT5TSKmwOe+jiDOx8jzBcNe4KzGrw3rBeqtJ8A
ZsxzAdltJr2uaKBK/CzLqwaPgT7DvXlBfzqbKNXm90W18ZZt4LLgbifPCZvaqxOI
tNQWMh5g3lG9ZTr5sKFHhp3KfoURaLX/+VqgEXMJs0BBFhPmwusfFdSqSF9p57Rd
qVKS+jdEYYWy0ecyMc3/P1JeuVhrTtVVC7cVsBaGLXNv7gQAOkEJqRRXFQKJE5Fg
OBSXzWKaRDJKAJ+R13feslgvvdNRzNWlAEEC1yRS0BR37qMMcm8W35v0pXZPJNKo
HwA9typhc1OxbYX1KI6ymqyW6wYiKxzP0VKeprYd53LI91JQU9v7RGYh4ZMZWPdM
qcdmDpNeIIcEfKjHplPu5VvDXOxPSHKeTaG9f51lojfXJZVGYfisC20DYGRDf6O3
29AoZJGEvcDThs7Lr19EQRGWi/7gdAvHGuMFL8WywtwY+HzYwvAG2AbwQKKZk08a
IjUPTkK4XieixlPjoTqtQx1V4kkhCCUNEhXs/STgNMVe9CtEmgLdNVtLLWGWFP+8
lCy8EjWvyA0gPiYekUXa+3g1iMIP0Ncm8JP0qPzQ94suWs/4HsYfDQz04K8Db3Be
gJcRyCmJt6mUQaVFVVwr9bsT/kpF2kyX3aZ7GLA7xy0pYivC2VBOESWps5DAdvpk
fV9luUfVhNRi5tDeN4C0aYOV6DIUnH49KshpLou55CgO+2jbg/wZVrJC8jZDfMPi
WPX8lqQJoM/IVkKpwxCgEPNiMQNGHW/jmg+BKfPoH1SrTNMo5oXcnwJufgm+pgh6
2F8kCq/EbLaB4RYMbhV/7cPVEOXrlxUhK9jKzZwZyCoutW0/d1epg2Y7LBV1zypC
1DsAAbMdtThIzncisXH30Mr4/swsRmyBtb1o5kVEGCm1miq7l8TZ8xOalaMK5O4R
+X+/qbM5cLiCEjgXoqUcxyt9reIlBwyK6aRGtLoSzIKMnkCITnqo3hcWsuLxC+8B
iA4OiSaVWi8BQBhL5bLGHF1UrN9mEbbQhY3mVRfmgV0p7HM5dLRes0llSS0qdSbq
ndZrLfdWh6/oI49dxN3tsIv9BKjwGBmHABN7m+j7PFducC8s0AVlJ94UXp8FMPdf
ebnMIrQjXbptvm2yDFbSQZ770/XmwIsDTxGzWWwTVPS78cx2iJ9hdsmek4CHI+ZI
u5xGDR9lJ4j7VOFwykdwIe0wj3nuJZvzUAA9IfE3rLEs49LpDaQCWu8RV+Yuk31h
0xe87nnEQSW0Ir8f2J+jC7DbUJdwrxvCSG4OrOUPJaErxsbaV1JggiFlUnHBoRqh
Q5dzZjnPLfxXv1FO/T9rRR00RoSemADw9bBCbLJVdluSL+VQKUntcWpkYn8eFhBo
QTd09WCTuh99M6KnVG/MH4jKVG0aguHALCTMYcT5p9xIen/pjEkvmqN8M0pogVSJ
qsJU+g+sKAZa3NU6udvxJCoi/HJatlYTQFS8r1TlwlsRpgQ/yQECF3dUawhdQHCy
OEirrxqqqU5u2rX6HeZRgDaONUnZN35Xl+5BqA2PmAXV5lS3I59gSTMyQVgHEtRn
NQiB3ysRTosSM/bAm+54uCZa74Q7LEKUA81j+5Qaj0VlMcSW60BrD4I+z6OKIMp6
S96FR8lRovXITzGlEV9qLuvwOcoBGoPj5DJnSfzfKzBONAsfTw8lEMTB1Elba3yZ
zAzQfgbEAFtXucaF24UAL9lmiOT401HqVw80Hef5rpQzrojqRDcn3dPrY5WrMBOz
4l7MAqCr+MS6YeBP+CmbyeprVG8q9mbm3cmG+o3efaDb/pTFuC21jGPTlJ+duu35
ycxnWpLX6BrqL6OkZlOQKv+k/WomRBOZcLOi3eeL02cs3S0m4zI5sa3Ak/Dr6wVg
ZHfUcXH4L5OLlx8RvZnuvIkUZSBwMOfoz/MgGYaSc1LChKRlL3iLdp4K5hwalqR+
l+QApma4baqsyglXRKXoV0zdKbvudvwvn+A0DWOtTFWs+jrYqyJm76WmXfNxvZAk
3Fp1KoCvlL76BcJIcpD7QSkQeIJdDcu99Fy9G8PbVb6+mDJCEmt3K0B8poiqFrEJ
gD23vYwuMKHQWGj8+xf/8YLuBQHBHm0f4JzQBD+lcVEdomaZh5L4liHr14OrV/ON
g5xcKHHKfDMTmi21PPxbISVN2a7at2xUgKXiwVEJReM/gpKS1ClKWJYhoc9iqrEm
tAJYvQsYctn67v0nY1Hv+Ke8vMLEXXSzTH9cbw5uDpkULLlKMn3UpNJG9VVe4XHw
6YM2ZpE+fJTWSCbo7Yxgt4KlIEpK4Wnp6rg9AISCjOSMLZQN4180Jd2VGAqD7xcY

`pragma protect end_protected
endmodule



module SB_RAM2048x2 (RDATA, RCLK, RCLKE, RE, RADDR, WCLK, WCLKE, WE, WADDR, WDATA);
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Lattice Semiconductor Corporation"
`pragma protect author_info="Lattice Semiconductor Corporation"
`pragma protect encrypt_agent="Radiant encrypt_hdl"
`pragma protect encrypt_agent_info="Radiant encrypt_hdl Version 1.0"

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP15_1"
`pragma protect key_method="rsa"
`pragma protect key_block
nasInzj1iuOY58I7LzYgCzfJ84yP42rC8jo/TCXbXNG4S9beKrj3jtjGJxahq31j
xdj1+v8iDZi4fttEaOxumOJhRRhIl7QxoTTrW57AI7Op50qHhvwVzcS7/IvYI4hg
kwUP2If72enMsoEa0RcOEI6i2VSHIU3T3ZxDbf+gAb3SqQY98qiiRJobkfD2w/RL
H75NZ0P5OIdIgk+JdbdxjQXhusmjYKtKDD8zlUhVBkhDlUSE4DWZTEqse5J0pqrk
0sVd2aSxLc0lCuyU7wh18yjIUkBZzLdqZ1u/pvUVDkEnunCXWktWIq48ijcRl87K
zFJCLpwE6RmVZTXISTOCdw==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
ck6ISNGVFkiV7GisUwb1C8vS0qFiL8y1eTAoFw3N3owbERahtLt+FnMa0iqzYwz9
Qlq2gMUEEO2LrwiiZd/GKiiy5HilHUu/L8UM8ja8j2SwAsGcSb/MBq5WdyJRCp3l
v9ztlNxiJDviw6i2E3npzz7wQVvvVoepNDLIVOqxFAD6xLkHxnlGfRPHMLqZEtqj
+S2Yb5mykEGe8wAR0BphACY/gq9AHgxtUHWi50UsXUiDDsNudSUQTtzflfK9wTDx
Tb3sXA1UxnS6mrNW2hfeX5lCTNEFhNYXnkKq86HCZ5Ng32QivI7L5tAzhTkqEfuB
fv+UzkkaFkxRvebeyDZcpg==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-2"
`pragma protect key_method="rsa"
`pragma protect key_block
NU+SIhIh7xzqZCh0tkoNejq8CAbDlxbbUCS/aFf2ZGuY/pfv/Zi1bT47ok/L0441
jmI9PopDNrk/Z9jMe+Xe/CSkWcLTThs0AWE8uxek9K244snS6uWmM0LkE0VciLpL
RXfvI+j2mL1YVduaUd2nUbIK3sIsWnjHJYbj9lNnhfTPPB45YH3KO/kk2/kcd3it
sHPcjQ5hapwkjfMHEc0Uou0UnJ51mHGUXh5Lb3rHeONkzIp4VShpfz2sr6xH6a26
IZJSO21BGPwuyVzg5uDUEYsZ21GL72Q7Feww7RRNznoBJAdtxPemCwdvJPlZBK7x
jm9833DTE5Zf23PNMxGJfg==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=128)
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect key_block
aJVetEsWfLe6Lvk5BQkHd26kPGoEL4fsrdWbmJQWu//7kbs4TwlHi1E29eHlU0Td
9RBOIBwmUmMTtfmKtb3ADg8G2ewQx3MMIRVFtqGoMAUGxyBXnBxqwATch/cEFTNb
wndX5Tk0VWSyFYZTEQ+n6NKhYB0wvcyWfBOlpxIShQg=

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Aldec"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect key_method="rsa"
`pragma protect key_block
GqxDhMnPNVOnd8pfkZrseQNxyLusKlB9Hc+2ht8kNsckdFoBu5mku9Rw75xPHf9z
APKErlvxhk7+T/2OAgEA9Qdi7E8Zk9X3lqAuzzQkoHFWyEUKnQo789BqkxGL5Q0n
biKCJFMnw4uuN9u8KoQOO0wZ3YBYfCRPswbEn6j9tpSgT0QKroMkyG4NkCXBes5I
a5XhTKnZxD2tMBVakKBvhTgscgawTMZykKsu5Hz+NU2IXcTIdLBl69/ZdrINBxO+
nKR6KbR4Lu+XjYXsvmHbLzoptcdtaRbHXJgmzg1bLHmBASW3+4c/hcr68gHJL7cp
CF108jLXE7t64ic4dEBw5A==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect key_method="rsa"
`pragma protect key_block
k8pDh7InTfyTqzvAyE+iaBFiOfALmWHyFd9w+zZ+QoC8+YeyQthuaRHO5zZRIHGy
gpM6B7g2GEIjp+8+ggHokmf8Sz74FEGItwmIvbE7NKvSdFUYRL/gu3NqFZ1UPJMA
oriTr+0C/iUOmT36Yyzd9LjByipXJCOoodM48EVO+ii+jAi/wjWuiXOEvw7zWdV3
vFCWl1VykU50++YlZi3zegNDvqPcNwnapc/STpWaqcqGWPENn8eMQ9tGBsGQMFHP
RLUzp37Wk7sai9dyRCh7SdZzXqL3K7ifx0Y8tY+nD2LgwmUjXl51QxlY9/lbR2nE
vZBuTnGLobXDJtPa6XqQbQ==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Lattice Semiconductor"
`pragma protect key_keyname="LSCC_RADIANT_1"
`pragma protect key_method="rsa"
`pragma protect key_block
V49QgLuquzuugF3+08KbblbXlnn+DDNUtCLIS31OfpPiVVN2mOKZsq+Vv+WRvjMN
JZm3c4RpGWatHoPHAu2RTbUY846tmnBmwyytDZd2tCxOxSahaLw7X+mwfpfluX+V
NT+11FoPszetUIpWj17CfKnHr3OIXOofaLlZSdl0agD7zV5I4MPxVhzP5uPKB7Ed
FMdYEHoxPENwJrD3ZyM/f2h2lfvwdJBFiL/2l4bk2hP9IzMUb+x0w3NMjdzN4ZD8
k2KFPk8e/piTIh6ueptymLUU3cuggEBAeEVO9XAK/KBNE8eu5uR6CBm5T6EkNtCL
KhwHoaSQIimle1nDp9tSjQ==

`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype="base64", line_length=64, bytes=3856)
`pragma protect data_block
sXteoIgnIrslP+AbN5py6pN7GqVJVUCS7JboNkB9f1t9Gk+FKrResavA7OBznXVu
jAO5B8mD/edy6XIjq8++s64n4juP7+bwN3OY7/uzdxsFkix3H8911RZWszIcf3m6
P3px/zx3vjeLXtaqBEy4VnEdvR23Cp5n3Vex3uO2c8BmgXcs9eBQycE95V6ZfCyv
d7752RYyg1hc6uBVPetDZDPSkI3dise3X3L2pjKpNDabWPYFI2kk7/Pay06EnzDA
OsNUKc/tcyFQeR1IuibvcWvr1i3YP3mQ7JF2E9N6bJ0Fpe/EmkVRf92PBvb11mON
lh8NQfexUiAxrqi+3mnErtJjyGzCTy9ITf6u0JmSPpgdYh/wzbxi+BzwaSKikzof
DEUjcTs0kMIxnTCilt4hW8sOdmTkcQ+c8PUFTJoL6OktPqqlN5kJ6fdDqDevo0SV
a06yrE0wUqN6NcEpBYsVWqqQOCeVYRqYhj++uG9hAHpghjqBcLHzEKOzIKGFg8LP
z2oghShlsk8riw4qevAiIOUr2bLOuTeTzskHzT5h+15wcYsUOhJohJ1NxwKRlEsp
klkA5tclG6IyqlRXfLAAM3sF8q0detJKlCxFkBZYYXLwyIC4P1/iXG/U/dpCjG1E
cn62lRIfnO3SUdvf14inBmii5KanRz4GepcMRXHb7RjeRFrLP1cVKIOINBmj4ill
H6FCsvXc0F6f7shITx6kFvSOAgnM4wXlSJzVaMCgsRKMMsoAQyDVhnSG+3cknFn0
Uhy9FtDFyDe/Ds7elXts72m9Wu9DdJC3/NuH0yDY0nSuR31wjtik02VQPmH9rPOS
UGqDh9DAQNXjxWdX3YZVvIdRc3gB8rS77zx7LBtxkE9yTDxcmaqZjzxLAQ/GrBnF
DAjdKBXWB1/UT372OL2G/LdOX0vfw5Z5/NavDcdcK9snEwwpkfasn1yqicW6Ltyg
+M1MVQ95m/HPT5A4h7JrrUxLtqYedx2aicuS05DmH2saJt9Y9Jke5/E+ZabGYx+l
q2zZMg+/Ltjy+vmDd6Wm2W5BPAgEo2SXK4BJNY1xdkKbtPkA9F3LOB73HBmezcNh
N1sbqTYKICxkYFEUula1TZH6toEBBeic/02xYo9GA1TsQ2Qkb/3bKearArcT4jjg
ApXsi1nfbdIuA8S8t+tst1fhdhkyL8NBy9VDmbweUc2ygtB5vBz67Ou+3W8lQyNI
ElibjwYRsHUhYD4P0IULiKynKbld76y7udybOVHVayPVC+BaUWdIQHUTvdNQavGC
dNGYJKA0nGvFMVMk7Tb38OlDQZ3/8Rvjxj1q6MmOQoKl0FrGTio/VylQo2uSkNOn
Zus3MejNgU21NNRvvOynZ79ruV9apSE3LW4dwL/eQlP0ubXkLRFOlqjNBaEkLTl1
5Y+/eDcAdh0s8g1SFj+5e4t1iMdP4L2u6xEe9A6yU3+GBg4O2ErY5ZnlTRUBkLdE
4Hs6PPGCSAsLdeR3BjiDKc16HN9Cg4iT3qrk+jQdZyM2da4+zls3lU9oMwh+v2jK
fpyYElzjo3vPVQKMS/qusAlWZF8YW/YaCZfiWVlkNMUa3q/ccBluIhDbUvSmbefS
Oa1WDhm/u5EovOB4YjBvL8XxrlMIKnJystQbXz9kdV8AZYk/0FD1oUuM3UfIdnzN
nDxRidmR+6P9U4Jw9NknM/ZGUGHh2UZsrG5bBqT18C7DbmCmqMNek4cPr9RzSO64
wKdPUhO5gckZvZebkj2oBsH+Le+/2cObblY4kFtz0voHwPdz60xS9zshPxhBeCBH
T8ntkY73B9sIhwL/mYpnFyAOUWsbnuh7BZcmYg/spWvPdB1Jx+yKBD4xgGEhyf0y
qzTl4+5y/v5RJN8K5+/rtgUTW/r9hLCt7wWGT38JtA+hSHywSNvpgJJwtl6vbiqf
AYv32fPqk52AA16EKNCgoVp6cvQTSVepMNjHEpAFKVoMV6zJIkiXhWja9mhKwt3m
9G7TmaAtkrrTy08rQdR5B7Iqt6hIhIKONZBgkO8IgL2xapMjhKYJGqvKpcLhomgw
G/VJKozFCjhdXUREZKDQNaMUq0Cz2YhGfPpvBNvolEA/EGrhxbX8nt236UHae9mc
WWo/lc0S1s3QMSYts5T2XGL7QB1CKj8PwDvBKyhMl3QibhC3SgCT1qqLQu6hnkIE
lj6QXs42x9a66bolLsbwni7aFylOlJUChf9xj4mOMWAWzR2yecg2QAfFtzEgS119
yb+V8N27p0SswmDZW7fgVh67obhOrSe2beBPzZJP/TK/tnOYYyGiuKl5yibLMXmw
2jQ8AKuMTBhU1bNPAH9trymJ+PK848BlaytZZkoi9yD9NB7k4tElayagU5iKxn7S
MiSmzs5OFFaPOp5Bq07K0wwM/4gR5w7/QOduh7DdH/OdsOURgBOCtKJ3pqIkyVN0
f9bDPo5yu2D0Lf+GfHCkzUS/qNyvoPvhqXyGwD7nF86vWrg8RgF6IffLb8RBZ+qh
X78Q33SnJ1oSlS89F8HksXm5XRKC0Pc8UFy0u6H1TstFsgex7HY5AFDXb9KJ2HPx
DljLBFq8cpsFq1BrQKEGL3NgO32NU5BjJ8hqQ1Fd/WvnmjQt79H9i60f/JG/c30O
2vX29C4ORejcNM7LFk+IQk3T9fdcP1oAJyAugBhWCZZuU/pNWVcpC9nIT3Jb8uew
7mqwamm9qhBp9YJuoYbv4iQ86L/XbD7CALINyUUnu1XPWOFFo3kqBtD0IjXOXUrN
ORr3+D2kiwK9nl7xEtvNALXkEVgMDgu7H5oLtUb1dDRm38M7vdbc+FsJxGqZg4NF
Dm2jywZwdwcq4+TZA65rNBJbjZErK2MHvGukyRhMgfd4hxIToN3VWef87yk7MyhE
Rap1mq5TbK7Jq/fcQjVNk33bO9cpBeE1Yy3CauPdq3aCwSe/rnM9vUYUv/TN7OCm
FfR/Ds6Jk9jhsV5UHxhQswcayssHOpQwPrfeugwE/m+85yEL1ZZPSLX5GW9TY5Cf
Zfvo1EK63IHh8W2qJvBFc7ur/kjHNhEuXlgJRTwIxROAIbhCN7jWHnHT8OkzFE/c
dvgz3xTMFFnsQAERHxr+FotHW/8sa289WvCJD9/kKvYmofP/CcLH10f+uzKSIuNX
zDzu4b9aMmEq0wkseE2Brxt6JC2xLjY1cJgFZouXP/YiuxOhsi6X1+5b3joj1Sh9
4lftWvOlpo9XzN3Q9CmG2GZcQbY3lNVo1QtBt81nDEvXffB36BC7+AIFMTjLzidx
+JtTtxsWiVyOaWXlUSi4m8rylN6E8C4Rp9ZwxJHB9vzPsi6oMg+Kwrr/wFh7d5Mc
T68TTsMVlS2Yi6KhDGZB+H/Bw8ykPPA+DRZUHTEheZNY9+LCgV395+FFxg9yyPBt
2aqhAQlGD5mHYQ1kVSMwdSjIFHJnbZnV6FDHX6aHseTr7rOsmoa7AVnk7xZCIadh
Tmfa/N8DXwoXbZbhkND9n3dtwMu8sRnlJ51FsLP1capO+qUXqcbMiYqXec1c128R
652jloNPGSYg/pwo+mTnTj9iMX/d0uppKUbD1eEZTP2KxNnrS4WSQTFdVCpoHOBY
ZRjNTQ85NXQC3NHZs2F+Q1gvVJIr4NcsvY66UtsDIhUszT5aahJoNSsAD3qDHsYg
YlcR16Gu9XDiMCpDj5M0LykPzrQaYNo2vQ6StEklZNmdPif9icpvXUGV3g6tTTSu
y4TmyyzYqcnyxOAbXWEi2vM3aKVoL7QX/xuD6VyhgrgWwToEQWrZ6etepWYphl5p
ooWy6Z7GqOct0Odeu/eJhKRRyjiPTwxloLY0mzXI95OpmziK37HqbGuB6mKWxWBy
wY3Zok+Q42zWE8jVRSj0KYI9CHyyXztiJh6A/27ACqUhfLfVnFuPGWseuYvkkcUS
LrYK4kd6rFDi5GfjOxL1lCSf2bLkKGB+4juNMHFTjFUUBefzSlYjJFyWxUN652j4
2eAbkAp6rF6F5ds/huG3rzmk4VQVUBiXmoa5wOwhggFFAUWUrLyY2ZQbgQBC0LIZ
Msb8F/gO+rcigV14eDAHIShpT1c65qim1NBnFbLbUcmry3QCjU99+AgWg7CozU3p
wZYk3+CfseswrKAxnkQlxovMoklbOqd0+b9XclD3UCQBX8DUkhU44ya/1mqt0gXw
ZiNhaWEw5db2lWKOn6vCahxh7ENxs1J7v3n0+nrgxlWlPkfDaa0JadDwGDOPImyG
H8zLT+yk5E5F8n3EfjrT76f97/xxVq2tGzsAFsBGhFGgavjjN5VodU24jkwvxuZe
2MUNptXkTJiXGKh+GuJrotHw08kpdA1xEZ0jmE9f7/8Jc0HSrRec6s5ZCscdK3HO
NLSnoU1N7tOKAZMih7jH4uVSBLj/ziazEa6IHev2QdgmGdA7gngVewyoEFYJKCJ7
wFTk+B5KvKGeS9POLBEcFp4hQBopTQoL4NCDrjLzbcsyYKsmzIxfPJZCAcCTDG+t
uCGzq6O2AlIwv/yHh2NY9MHVgx25LSjPYBNFnV13mdMrxpyifUrqpjkr+Z4UO8a6
aAe0cX5yqSO73F+4HjbNP1UlBYf2TdCvCifQBV1A1iX2knyghr/+fGUKNdSJ24pX
L8FyeI20oG34mVL4QRF+0JhnO1cKV1lb1JKMl6ex7Qy/yXm+HlbapcoCcXekc3fd
S8czPW/Vib4qoeCmukyDS+2ecgFg8yYXn+GJU2ER1+yx28gVrO7RzpZBRQe7S1b8
L7iPN/8LMjG2jKix4Xwtv9VJQpl+6AR46IU8nXEzY7QdZFRHYAchTV9HRCcBN6O6
mVvReCMIpcZEz9HcAXwXQNpqE7rv1A9Z5pkeEgSNUB8gXva2vy4r/2mqMDBUAK4v
NoC6ODHVta6G+trtA171yFlyxQoLbkWLf2URRLZxLVfqslVb6tlxN794P6M7DwGK
ePTECGtZfw83u486PhWMCkZcIEtV+PHz+2gxz1+AJ8wnQLEOpMsKvakTIiaaR8mQ
CTRXks53tM7uGwJfLlem2p0zkKfiTStnFEOdBXbhMGvtyuvKUBsP/9GIJZLwuDoo
d6LEX7dBIws/sB0abIjp8YBPj3fRqoQiTyDFXcFkEqvryrQGS8jaYjQ6tZpLnIxI
eMPc7+BTaWpP5Cb8cbTjWA==

`pragma protect end_protected
endmodule



module SB_RAM256x16NRNW (RDATA, RCLKN, RCLKE, RE, RADDR, WCLKN, WCLKE, WE, WADDR, MASK, WDATA);
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Lattice Semiconductor Corporation"
`pragma protect author_info="Lattice Semiconductor Corporation"
`pragma protect encrypt_agent="Radiant encrypt_hdl"
`pragma protect encrypt_agent_info="Radiant encrypt_hdl Version 1.0"

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP15_1"
`pragma protect key_method="rsa"
`pragma protect key_block
cZM9tsBZ1yyaqOB+XcsmjmvWYz+Xm5pLlBN0jzzh/b3I9z7JR9aDPsyUfyERNnIl
oybN2/GDl5WalwEzwWWIRSWLeJxJdXHshm8lFXDpRTxbz3deFFgW5eV2NTwk3wkB
1ZCC6/yScCPYXXdrKD0QIdNp2S2ieGvxHNFMUDHUJFO+e053DjXk1oVkDXu6gGsz
EvWdaRoyT9BItTqzce39GuPZEgqHhJppyD1X2lg9xSia+efEVPRYpNknMY2TbMrg
Ge6Uajs+ZTaWUyN9TsK+4mlpHZ4LRRA0nKEHsNHpV2xvZAl3UaYTYI6vyVEcVtC2
kblvzcygJFBPbC7LlUb9Tw==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
Wzhp1awJpI5rNajH9yQr6gC+IQnB1SUrTmeOR49I/biW/Y7YDYKC+7oe5SXL8+ZK
t2RUF+lMMmdg/78jg92ofSyfiQAIbxz0t23qq5Jh1t1eM2qf0IRVKv+ZQA3MKhxj
NQdD7qpIW5mC5iyXk9ZwSxMdaCBOnLbFdpvrL1Gi2a5oJxo7X57N9+FtFm9Pp+PY
lsiBFNH+B74M1qB6OEJsPMxv8JmnwRzkxfDAoCDBIfUnYCQtGNzu/cW0zNs2yyIX
hzdrzCBDRwmIo/hSO1Xn0RUMxbumSN6UO/GNnKr+vVKZSnH/LY1zSrsZk8WohnJZ
0a8k7+KY4dkfuSD6fyQe/g==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-2"
`pragma protect key_method="rsa"
`pragma protect key_block
A5jdxRyTkOdz8/scVI9WEqJhrZVgfkOVYZY3FafEzFO0J66h1Rw7GnkVu3pNuyNy
6Qo6CFv9k4IOuML3765YYqAVBTcc3c85q4wV+Hl5ccFIPgyjhLF1mJNPJxpSzfrY
GK/lFV/tO2VMPmwKQ5tnJSJ6ru7P9qTpsdIIWUfkOCzXSqXbc5YRyWaPybhrZlpZ
kPyGnSgvJhuc+99ru+Oor4trUjL2DLVY8RLKs9haXpgqNcDHXLflIKvJuOkS/iEs
XCZAAsEzZtzfnyLFwz3BcPIdz350TFTJcCQG6BJbbBzKVsndBeDPlTKQjz6rb0wc
4V0FXjv1/aSJLVP7gOMXPw==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=128)
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect key_block
ynRdm8iwN4FcdVdI8X4Ch/pygbjYV/KRzjE2OhNk2USAB7PG+IQkifzioo2iU7PD
ABGqf5D4DnI8c+nKlM+gTmstUgdxm1o7zX8Fc5mQ/20WsALKS6Q451Dk0rgMDiYt
tNn7+C0iR+XIwPoj5EgdtitowA4TuGemY5kJM7STdhM=

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Aldec"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect key_method="rsa"
`pragma protect key_block
LvgHmelZ4twj5xURX5H+3h3j4U+v2etXNd3n6T2Ax6ZCW9zauQ9opgSLvBc7/gzF
W3cNGB1vB8QdmmtBLGZHScENdP0o1XrcKjmq2vTN4tkFtYCwnm6cWQ5wS4Xtbush
1sLmRqYI34mN9MHxR8fbGDzKh0Caoeb+apLbWqxndoV6hqkXY9fmGw9bdPaF3pPA
joNCa/FCyjlpMHmw/8Zs5hoy6tM4ambib48ADzxJgUkXcGcPAVgOv1cowrA6qzLY
3kPfPxPJIq7KzTnh4KZy2KoKPkku3BWz5UElZjPe493d4S/wN1uMA6HpkPicyWun
wpEAKnyRAwysIso78ZkZqw==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect key_method="rsa"
`pragma protect key_block
IZxVW/9GhFZQMRMMfNve5IGQ1dOPIHPJzbUXTLWosXHftrZNC7Bx0u2JXhTGRUN0
qpwhHlecbUsUV9caMz80Q7R9W+ErIgkm6n5z01AYdwxpLB2mRSGl35fHUi/GO5bq
V4k856A/z5Si5ImozOOIM+/nC5Plv770Cn1DQHljQy/T/3x8u8cP0ERw2S32BqvB
IOFk1BOUOt2g8nwulzhTTmIYHpRTJi2xsmo1NEfzSQCmeLT25HcSz4VxJpAlf/fh
TERru9gfcx6vOhv1LP0fi0KbubkfUFy1sXsZ5jdWMlwaFKuIC8GzgcHEoKbC4aYN
mJOgKOU0VeuAcuSl2WQFmA==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Lattice Semiconductor"
`pragma protect key_keyname="LSCC_RADIANT_1"
`pragma protect key_method="rsa"
`pragma protect key_block
pqmnLysPjw0SZSrpNnafUpAF8/tt0sQUy+wXIZntzN3k/3ySkiaVGmlBE1YlLxdb
6p7Y4zyOJESBWX+wOpEqvWaVuUK8Qk+d8yks0Vg9ay4vZ8MtgDVKPPsAhSJuZ6OF
FD+uobqOw0lB//R7KxDAWwBJSTYmZcfHcrDM4Ww/6CFRMRe17CTmXmM+cFARUNiE
6PGa16cnO1HsYsd3yt2oIenNcxiK1uT5SuZhnV2sRXET727kvgAEKalEHs8CQ5iU
+xkavxeotJkee/N6d31DdSPhqcSt8tgROWOJ529MffkG/1knlilvSF/qycDlqiP+
cCVb5Yb5WT1aKW3qb/BLlw==

`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype="base64", line_length=64, bytes=4048)
`pragma protect data_block
kliY0iV3T7hIxJi6bXaRwdNCQwO7+8I7UvkZydsVXPfiyQKC2QhCP55bw0TLAFbF
IhyhJT7J16CHeOVEqJxS9STVI3Gj1172mQXYpspy0ed7utdCxVLyM86MQSwjM64h
YeZKkb2Qqn0gvsmHynwRwirbk+jI/1sFX6p8ZLmyOeQR8uuBwuwUv/RuS8j4t8KU
TcxYibsWHcUY/32Z2gwtrBGoMmAwD81GVolJCWmS7Hp/TC1wZ8jIqfTp0uZDDj2o
FKMx6tEQ12nFFfVK34m15C+6rtXBVEkuazSCb9vReiP5o0jam41RBmiqKlbBc/Y9
T8ij44LteSd0HTPapSX2ZVawI4+IpKJriQTReAn2+rqqL6R5sY8vfUnfqk8j1AXE
FbZ+oXWbiVvtqQeRHeTmifgX6IH3fCgjq/ds58ohVuT12EjKq3f4m5uqCMw5J70q
kYK4NE0BDMyxqT0jJHqDwoitzg0rbRcXR+WdldopEJKPuozZ2aSqKSTDJVvrcWaM
AzecE9RZnKMSa52TRD3a16ikWMr5ocGACeo9ZRjhdkOi2j4DGAMsRxeDjRiwQrB3
8mdGvlF6M+kOrYqBD0+CMLxN/5lwD/uWcJv/n7l0WnXV/zhLDFK3LB4ubxSfSFBX
uF0rGHrRovNwt4B9sgBcAuEc95jjJ5mVfiv2VUNvZ3OvxnAnWTliB+jXcjTcmHov
cOxciNfLVnCSGPW6Jf/6Tt4aNW5PppGWM69WVuKnNuxJNcyDfKNTcuP/npFNYUgh
Irmo9V0xwbLxF6/9Tp5oNE5wag10ZzQIbyDbHA1C6wBJzr26MsmXxAeiKReKAKlg
rdjxkbwq1P3ipiFjOab9l4so3kxv4YTM7EXl7ambkvfgkNwC/tmLGqcEydZY4MKP
QOp5n2oUwSrwLB73S5Pfgx3JvxscdK12MYiWZ8O6Oy6V42hocqQTZ/cE03mgAF0F
0VnQV5zbvEKk3PfU/79Iq6MHfgV4B2YaKSDBU6A96SGQqGt1odMIL+7bS7GFHFOl
2AR3TrUtd4ssCWkWKZ759kNeZGP+brA+d3mFFmUU+LBAJuG6nZUM2sZnMaFOq29b
HBmEyY8oza0iuRisbgPet9SFgKFtzh50z67kSg5mISgwG/0BJfKrtEG0DRBHN42n
kKE+uTOfBO3lI047Kt6+Zn6Qx8BCyv8Ka3dhPsVVYdrLxM7yarVuNr5JIIGkwK8k
rwmSefJUvHImqIyeSyvUteJwEzydH9vy8cS/LKBGklr1Qdc8r2QivOqYZtONuqr+
nc0IY8XVCEN/a+Y+SiNjsCCQqWPP2b06Vky6MZGeSvdgTBU+4UZXujUAK6IqoKEY
MDGFbTdMGOWL3mBOIRkRLSODTYNxb0tG/shoLamlQAYHUrF2J52h5XibVO0eimuD
mPxB/zIA5EXGYC+ZCJHaH8A/q5DdWIu/OX6jTc2nFvnjO/ESc81d6WjXfzQi411u
Vhj4B9mLy8Ijorzy2NDXLhRc+saQPD+XilAcTEIn5dkf6iTEcu28CAsXa4IdBcDt
blHdQdgK6cX4cEEN+bV1UdTbW1Ll0IOjZWPmvAKVvhe2AzP9c2xotCYOB5c5TaQT
mH5hVlTzmvduTmARlj5/0Y3NebvoNcIF+J3vK+4zAU4XOHHTmBqhgyXyGxNuD+dP
tCLwe6R2Tod5rxnpaQ7XyLYm4Ru3ALEbGM9XvNKkb3EQNiKV4uJkNx9EQdKujxNJ
QB1kCStB0cpAYmHpVxqe1ie6CerngczDdjaa/q5K/qaZo7eEhjkkRw1ppX2SRLsK
7gayEpWBQdICvmXocpZg5kblJgfawMUKAcl3VW5wbmaCl6f8yHRjiD8bkQE4G5Y7
PpQWhDyXGtzjgV6JdjrIOa3wmNwz3Zq46Z2zGny38p31bqD14vHZlqS+A/2pJEKU
wps/52bjMN+xzbnETrQR5zDEy8Oz1N4iIoMSL4d7LKuVi8oSbb3lZlEsRZApQfN7
4yCo9qT71YpLFRqgLaAeBrMYbJ6dzHVhP0KTIjTSyDLNp8A30vk0gGXbhhoP5CF5
xxq5CtoGiZi+NTK70VB0vxOQMc2IS6+TQEbI2HJVtQjITvd8+zrO7fqsFw929tHg
vUmAz/EA3Uthgdpdvu8B/ojRxZeUjVZzHA28hrIEc5DCZ2s/pK83H/AAnsMlyV6c
QcPLnOko2X67/uDAdfzqTswJCP/OKHZePTeMOw6FrP2y0ib4mmrVLY9QrCYurV5R
muP2RMyz0DrQ26ZDys0Coc8EFr8HqAczRWrSshmYpCo6mR1ivfrH2jpkYRHRC2Bl
8q43lknijx8h2f6MhxFzLcJacMCXrueOc+3fUJyQ8hyv2iv9jGP0/MarN0tfSX9T
AXIbGZZvqgnA2nmvzogEvOQvOekgXXhLrFqW5dXG1Ul2WbZe6PGcw87ejCFnuX2T
mADRce4OVIYvMym3v2n4MoHINlfuSVq0snJit8GTMIDlqiwTT52FGWzqlEIaoe4p
g+b2blLAObzOm5k01nImySYeWHmVDaV/Dd5Jhncu1Ipf5e9rs8MU1mbz7Yc/TAr7
OVUHph9+1EJByLqAIroLwhkm85aTY9XRChhX2Tzn0GWIQZg1TAYqZM6vc0LHepnk
+WMjnF76b+3s6aR/YMQp19Hdclw2148IIYiD65G4PmWiypAwfRDl9H83Ql9XMSqh
4HNzs6PGcVXbdWXaZy4ii/xfzOhMuNWjfauGGqFWVQWrdnRTsbZx8CiQhoPZuhzS
2accDByT0SsVze+ehQMylDxcJ65N0tDxyY0NX3yQ/VXB+R071oe7V97j7SDza5dW
Bdoxt0VAouXd+nCljEOGLbH3jM1uFvpbdZ2yIKzE0kOomuVe7FLcTalis8EbenZU
r+CJztqZ5OyW61RPpwBlF+9uwBqF7WeD8ETynk8JBTp8XFq/YQEUWI+rIxBTMO7u
Q28GG0OomSbUShMuu1RdgJphZoAmrTCRmEDQQz6eUtXM3ayzZ4yky8vbC2aQWWyV
5Q9i4R2E4NRMlNH2WlgRLrGVUXQvAJjo6QW60rQAteTo9UKghNEQ5Hw+mVeOe3Yo
fCAjtMZ3cFcH6jwAflrDPyeb83DEoORoKcAmP7yrTTWHC907fjZt0U4xENHFHTZM
rGGt7b28e5WzNuh9FvvXYSjMlU944B+cBFDVTxhIOj3QCYJmw/c7EVe16RvdcKAx
iY8bhFlMpRhNq9xMKP445H/WoFZW9Q29FCqH58/NjEWgN1S+67FXwNX2niwVRZ6H
Qt/cP8U0QTtZ/EJC8pO4dBxxD2kvPfV7rso5lTh49XDwud3/HRWODrJvNK+PfeZi
mj0R90ASXdF5Ua7VeeZFObLmT2WbySvzHkilBXsuewOkYWjYr4ofwP3ty+duJi9l
AA+kshnvnVb/ctdipyoqXgftXpsr7ugBmWvzy94Tw6EcoyvqrmkqSIsjsK17mpg4
jCLgKhBK3uUbDsTUgMJlqtC6a3y5rGGYkjILC2iP0urZFHxtiXcCBlsG008BkuDm
pbTlKZZOPrYxjfYSsLLWaZbv+esw1hlMyy6oC456RmLix9LlP50b3f0JxRBXfuog
8wu2pYpHBZp8myAUGspbrzfOArrALU9fOGxuNjTqpDPbTKI5xJZDsFue+3CGrtdR
ihCbmhtLKpa0CgY90UCFTRa9P4OlNB1WVrWdb7uxvBL9HjKSl3UtQcTMHPJ92vvR
GVRSRJ09LpC++wWAOIP1+o2bov33rQ09+GtcPSYejJOn4YRr91fGkXdAi/JUN9/Z
mYjMUZgmCJp+miI6ZbVPnxf8Pt0ujC5wBVrF+m33987bBRoCdIkRXTFHNw7S4ag0
D4URXpj/10TV6D+QynDV++98nVTUYxHHkFW9Y3dxsx4Qj7Yk3e21i5TKLmhikYrN
6emIpNpJb0eByVNLMyHBambVyjDQjw6wSUYz6WAR8Dk5cuwJC8dcjGtm6DiZMYC9
Dy748A5kyYH9J7ssARJt76gunJoa+crF2zDi3cG8bycEQ+racvvy/h0QuytGr7YV
7gfFjcVi7gwE7Q4h7nM93Hld2kQJAP+rqOLfm+kcwWSjpQWHVqCFt6OsCEL3Xym0
8YnmOcjZOme66vMPfm5w2Bst0DnXwhO/mYGCaM2uvqIHXVwVPU+bjSun6lnfdU3a
TvWESvROsYnA8C8toN7Ci1tXxcn6fS90AzNthkh3oZXfmNP9ebEhr+erI/7RfK7j
xVkRzhtRIkHjIK4MsSpSeX2NGvuZN470BgjliPNHalSzkZCdk6NNrMGPKbh3vx6s
e/NWnu60gjD1jdBqXHDFMfNZXgPjibb9x9DoqV1q3LyrNnMflohEdWIakPTe5Cnr
6kSBRdyaBz0YBy5t+WwlJSKh99pIS/AbT2+z+8oU2g6JVzXasiYy2StRYaa3knWU
KSiRbqk+M3UXHA47xz7IeQlfy0m9n/9Yr9P9azlqA/WhMfKbqEnjpAXnT7/LOFgx
dpkSwLFUajEie6Wc/pG+6sZnd2Espi2v1R+T7JUolPJ9ePEajvuN0yf+XBnTbOqp
1DFJQ5I3wlRwv3YsBqEsMHh4IvOl3iukz3JjAHa/wqbxOpZuU+vakR4FnXBVW0l9
Izhp3wpQowhx9ZjDFlAYwDP1TgMMg0u989vUf45ybtieyJzmMYGUzMMUttn1EJ1h
TodA+giRaYZfxinYyicViwzXCOBpQ7fWUxe9/MFHrPIh9i99xTs4qlkvOWoRir4p
wAgrIc0YsdexW609zkW3+yqnTXOCL3MW9NEwXQjuM40/o1fBWoovczmkUhlcGq6C
8HTwxaL8zkcUZgGGFAdWqewlVMLmEZvidhM77HDjPL7OKwKNx7Y9ZBC87fRMV04+
Q4NSriGbCNPNJ6h2NH12kW4duJAZdcQiTlXMUEIcZD2JuK94yksCxVIhxVCHPmAW
pzFbM1AEpw4TXjCOlblpSWcwsk6gNqV1OIMhpJUtiBGG0WaWB0F3yMnKn25NE780
vuiSsyZwPdI5KuHrGDhn1XFWG8kAKc8/UC+5fEOtbmPi6eOCF1jo5R2N0Gn41OW0
qEP4uegtReoxohkCgsUGOBqvYnSgIlt2jikvPMubi9UIxRlZbahs/OTl+whkuy3y
SNFYwnWnfZvZOAjmHq5Ho3c0+SS6SxQN4JMkkIemLFQLaLv0/mg7iJnEXnk9UxTi
ORhOH43PO+L8AoVsrvm79kZoCylzQP3cSU7W7kifRxhImEErU3DlodalD1JbJSAf
qP6s1nETnQQeX1yrqkpdFeC4h/LCwCdyLwS+Pe4W3Kin1m7XSlBDQWWA3jH9/Aoe
B64+uYN2U89ZXe0Rdb2yFZyxZ2seSWaF3UnlKG9vgg6e3zZd68PqUz2XZgcmVzEF
6p1PP6Gl74VSUAvFJHxRhQ==

`pragma protect end_protected
endmodule



module SB_RAM256x16NR (RDATA, RCLKN, RCLKE, RE, RADDR, WCLK, WCLKE, WE, WADDR, MASK, WDATA);
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Lattice Semiconductor Corporation"
`pragma protect author_info="Lattice Semiconductor Corporation"
`pragma protect encrypt_agent="Radiant encrypt_hdl"
`pragma protect encrypt_agent_info="Radiant encrypt_hdl Version 1.0"

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP15_1"
`pragma protect key_method="rsa"
`pragma protect key_block
zv2Lf/e3o7ga1PaOP/P5yBK7aNJe0juZy7UhfiBTWFjTZJFRDAN2F4/nDFFIkYcK
aBlTRM9rN1Wr9yFJWInYX+raWvw0K+FDRLlUalmso/6XffJs5H9J7ovS8EKUEbKy
ZDdL8qOe5igeRM/Qdd+xftaOdMEnD14i0RaGJnF4fEDyL/22YmdWxl3WKQMmwJi1
AzbaVsKBptrS4U++V5Vh0Dy1vIUzNq3lxnHPiJFZyO15Ab259H0lAJ0SHjQ0EdN5
YDOpLTrMsVh+t1X7QPtXjuzPJdrLDJ2wxDF7AsIJYMygOeZAG8XzI43lDNqQHcpJ
Tc9fBpIDNzp7pBZILK/JGQ==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
aVcZidDo9+9p+BBRNHwg1x8HzzaChy0vkXWO1TBXcGWP3JXVA0lrL4e2pTKk0G2F
D437JayqxePkVcPfcJQo8Bf0tnf6QxX9g7KzhJsEfkOuSGuaFckLPzSB8Ft02ZKv
KNYoHfrvC1ZQfxY7lXde/vnSX0NBZSy2hfDIA88zHr69QFARNmFE99JytCIPhtZH
uqrQY24rCtyzQxx1fA/mVNoVgQ7XxGoG+Z4VuFVO5opsCzlTzPD2lQ1Q+goGkp6a
xL7KqIyTxVgVZENN9nVG9t1LQ6NPDL+GkJzMbNjQ8IOfphEfY5v9iExR20HSdmzl
XkO60Rfip6D4TJLSPipzqg==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-2"
`pragma protect key_method="rsa"
`pragma protect key_block
e486/MIpVVbidJ0TVcgTTzdT0tGSZB7EPbzd9kWxk5teKbvyCVCbdDIjjv0N4rpH
hn0Dmlxg54v+0tTMBscztI8jMTdvaG15uEt1Mt/jVZzfL2Uc3Qm7d5NXYwcVfcUg
hqHnfdVatz5wpb2GH0WRfZT9eT2B2uhX7nmeBY1kiZk4B4ON2YeAy0iHH3uDjH1x
TlmUnoM9cC8Mw6hTQxZRhFJVnJ72FCxsSq1Y8rH69x+qARKFFT52p8IVmXPX75nm
f+H2/5BkrtVyNeGwql/Z6uC22NCxYcVODrHdD+zEHzj6TzeRFUw6+u7iew/6UJKh
Rx64XfkwS2HLgi8gQtxXKg==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=128)
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect key_block
ELsrfuq6G0/FXtRb79MNFq+Xc7wV9U6E3dwq7Vm1sqb++XQoVX3hluTGkoQ5hh8v
sPYcNUI3EHEQjDtWvf4zaANAt57XIDGRtr/OAbeLYGezjem9I1uQkQuNl1a5r0Yk
mGRzIhgffw7fTzxumusdtxwOlYhLv7YHyU/17iFRFSA=

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Aldec"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect key_method="rsa"
`pragma protect key_block
owF1BoNJ/DNJW6UNZam1hQqCLKGD/6NekzS/2GIrfnyivwebkX2JjSwThAfTzbLV
m3bS/p1lFEHODeD/oQhdMwWymZs2QKPQGWK2urkVKx4vXMr7xIdX0CarJguTG2R/
MmF5YBOIXzxMyyX6aaevLTzJAe5faFta9J5SOgaQyTKABpCu6Dfeh+PFEBX5sbjH
qxYo3qAvVt5gpxcEMs7cd/oGpK9f2QyiM7BGGqgtpcEoEeMuLU978GGKPSULCH7d
YBzTXVzIKrZW1rFjS34/QY8+7BstHMbS60HwfefazaBHGR+QF1wxJKzbRnAIXLmd
IlyWNAuDJbHOhs8+afPItQ==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect key_method="rsa"
`pragma protect key_block
CyVTX5+ZeO2zNDChkdr2bcQ7/4Uhw8nVoMDkwYUdoZVOCXH1t/eMzzKyZfd2GEVV
D4+RPLDPjS7XOD/7WBTPz4px+/T8ns6IvEz9gEGIVADN3JSR0GKTOmgyg9rsjumi
Z8B/6RUtY39zF/UdNnx2jJ1NoVC82/lRi51qefg/aZ3GZS6Qviwupxaj18LwzFz4
gT8Z4NZhoTJav0JcgQZGStEBSQWs17b9Gv+uxwe21G6MpNb5yFEq/SCGEoKUznqW
LM2VaAIbFWbLUi3vvgDVA3l+ZJ/2WvJ+STAvQiz+Jff3y6vU3bbP+uKKza2ucfCa
RzY7oNC8r31WstizaS3HRw==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Lattice Semiconductor"
`pragma protect key_keyname="LSCC_RADIANT_1"
`pragma protect key_method="rsa"
`pragma protect key_block
etw0SEfvd2US+9uupx7dEEhCDILpZqPv17y+TPbjJh1ljggnob8xSIF1zBOjyhBR
eRoQLz8OOrF3R9EE8j9ZuqU0UkHXcQg8VBuPUiOQ5OfCPnIMje+0s7HJEk4g4+MT
tfI6K2AnCOWtA8BGygxhl1L5gn8yZ/lD7huSc4OAy3ZyqNKECc/oy7EKgu6C12l9
08MIPCOFnnmDlv0nIrtGM6ApaRoBBeJVbccc7EGk1TwRlHzjx0RYcYpKuc55gzVe
b1god4YCfEayYJWlphiL5kW/zQwp3J7nEGSGUqEPekQbPlCy4knwl3sbt4Ee7JN4
4wGyeiodxdcZN345Oz53ug==

`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype="base64", line_length=64, bytes=4000)
`pragma protect data_block
ybP87DgzwDRT5mMY6FQHKMSGsBvM41o8K2eF4gT4UG6S8TxhAIslidjypoWmnlow
tMRumXuFY7Cg/vyWACEwIQtlX+13BE3ihECJcPXNYj2e8Gfdc9IFrDCBmOGsYR+W
dGYPP1QOXP5MTmYLweCM6GYfDYJfcXVvfgv/fmSX1Y/CjQJA1HV1Kvtg35NGGRdC
aevCbzEiNEw8I9WSHg03ThsBwQaFdPvjDtcYRJoJdP2rwQRChe0lZeH7l9ALTM2e
3yxu4VL+NvFpn3Z9nsAAa0UYt0pdbNVYeUHieKbgkjFiuqdnptZBxSNYZ7C1Q8i/
fa5WGai8pxwyDt1C5IMqq0NkzJTb6mk6OuUyn+sc/vssf3IrwrX2MsUkWRvRHT1O
GM35RWlw5m2Jf6oX6NeudO2yZ/TI27XfCzgDlDxTxPvcX8wA8jRTUhki2BiBGiHD
hQorqx29xrxxSwPLrt+NyM9OGwzgwcBFJjBrEeWOK2JPR4s3zFe8gNMoMtI9wAHP
Zclw8UnV8OgTEwV1pxLeFjgaj2MVn0ftq8/vfw7cbDbl9P//YGigkzSGnAH5C60R
pHm54GTF7Zj885ZmF0p8ocaCSS4fAvp75z7HLcYgn6AC/wbVa9wSW0O3fAFsEr4j
Ow4DaAEvfGNU5FvaF2wlqS2I+NubE+3knlTOEfx2+ZJkN5p2/MEORzGPxIspipbj
Y0PtGn8Idr+P6zEqnEQXKw+blDLwlXL4Wh78548CQEJO29Je5+FouJKPiUofV9fC
SfNYQbZ/knivOe7I5Wtr2B6tRj7kDa8gH2rwLWPtIoGJtbZVqcCqkLnNu+0YIuzG
Vups3bPeu+yKrPQsIsRqeSDVZi9X78ICePUuK0fMbzYBROtxdLcvYb3WTQSmOY+z
dC0ZGfIC2lRhwcKU4KmKfZt0Ukkc/J0qfhGi1y8U8BEvKGHp4VgwdLWdw4/Bu6VV
7DhdMPmqp34/51u/DKOl1DkVUql161YlGeY19al+JfFXKCYd/32yZpyUXuD3vqZw
NVJcogPfdhMyFeDQZNkZoe19oGv956mmCb7EvTdincT20ZQMS+F78lhJ9sX97jjP
J8CGGSXFpC0BS280krQyryXKAQWLcDghDigZM+pZXIDfILdIS8QKNBlikapt0gjI
qH2qjUsmyXFxcdtOdsHtuiuzpJfUWYD6LTx9AeEBn6cElgYHYzHn5j6+lCRgiamH
MkpUCxlrnmGaHYFJYW5JWzrFGKmSUe7QUne0hAILwyKT3AyQGZgqyw3EwVb1RCAy
81WnDq64qAzXGWSUy55n0u8wMYEaXv8+xnH+ZaZIefft0HywSnKCtFV5pBNXDF+q
jlSD2K4fm3Fmas/BR6NSn8TPHWZjDcAs9glc0Srb4ooXJtdZch57KeQ4YyajKGyi
0DNU4kvyWx8D8u1Gy6IThh0ewo7JaDcKxv0c9lDWvx/r6j+kv2lsYGX951k18sFQ
Jr/Ln9yu89f4hzEkOevffce9UEcN/DPJ9On9Tmbq1SXpulNmOq7d1yT7XlzXNVMT
xubdfkfLETc6dgpyAjkbdet70YhvTr8aoDjtIx6BOz3V6ePgQKuXyqsW2IsNQ+rr
wv/1B6rlDyq2Fwf5pqBi8SnVOL2RH/zNQDrySiCJasL6LPTsONwQNEunRh+FdWYA
iLaPly83cHs0b6rrg3zOV4qtiPoO7V+tZAvEk16+7DRS8GX7cJZLCRbnILSDrY77
oRO0zOahWMPJjWYRtHzOklSwWU4rpXYHx21meayODBVS5JYSmUEl9EgNcP3RyKyf
I6wTn+oLFUbuR0N4Ry8zLj5q+D7FlUHTLAfLnolOinO8EqT4ITkd5QOW78B1CM6h
6fOGXTjhaf2+2GCS6OsK0/lFkxSssgzpvx8WGNYN4Bzgyss/ciDY5JrLMEXdxG9M
+W3XMHYU/uTIOifI++G7woyjoReGqGMEEiB4TLpY6GiAyutnPCO/5C5W3Z3ftE/+
uP3oHBGqU/GWmIYxBzy/+Tbe7zVGP31gdx4Yo7Ii9mEuMaOiHQYEE3YEnVVFQunI
2Itu3+LwIl8d0rFBmhyw3ISqM6/Zv/TH7R45ehfNErKJxB0r7lCEF583YadHroqO
yfJsTAMilQiAQMm58pZZsqq2xlvVNK9Ci68PdJI4kWjWnpXIzn799DGn5FtFjSkO
7tBqDHFHmr+B0a2aD7fHFcDJ/dGtpuPGrit87SzRIEXoTQAAwwgiLMTBQ7PWdBr6
mELP83EonZdYO9A+u0UpE8DJHGOTkPejLBn1pXQtmsdmA/cmXPWI+6nRvGRJiFH+
5Y0VqAzfN+SSxSAYOnPW4pobPw/inZhg1bTu32o4+JSp61SGTSlibccdHCOQNBqx
teV/meI/jxcr0yHV4rutjUe8ZA2MReMKu4ItPkyt+RUCb+89ZcoZCV+K9mj2Yiik
mMq2RPTNkGYKvnXvLhTOaYmP7bBREJLQUM4NVUZg9ukhwJ0xsLoCaKxXYUReRu2n
TeGi9bTfQPDTi9Idyv2HBGm0UghG+yQd7IrHdVnzRtS6lxg01gJggZQpG+RcqQx/
NQhgfArXysslraOrvZrN3sRytQ5xetemgZpzsa0DUKuIrTpD/01gKJg+Dc63kkLP
YV21Yty9RXqtgOco/zf2LG4QoxBNpKpDz599tV5mYMFzrPvp1iSqIrV0Z0HOaQzL
GXT/Oyfnzu2XTsufTsBxfC40iK2T2cfsKdFOQP3MSXlhloFdI5f2BY4wXTZqVZ4X
gw5e5Pv5SLHInfJ7HGHLaghCkF7YAf4h9KOmcEPdDdjLj5FCO3Uv5bvCndwAZTqf
4Huvl892PVeD8W/ILwnopUOKrsNROZYl9XOc9ZaEJWgt6SJqhJRhl++gBLvSX726
pCTBq9dBs3L2DUz9ms7z/wNdWE+UYE3RfMxfHc5/VVLTqf8lkY0Tp7pZhOOHqFKV
dGbgSOBqwxk/yjUev91NoUFe5Yhf9L8+AR5Roc+dQaNDzhyrYByx4SilfJuM4O+k
OLJQsv71SsNkkUCSMVIZt4aq34/zrhnSAzuoD/HnhRjCJQwjjlJawLYtQM8mhvRG
h29QtoyjgXDJwkQ0Fp7UhbO8p3M1qnDqx2yBvKQkU5SxkQEmfTNE58HFWR2Sh1dp
j/EXXG/9fk9KRKYikzA8pFxowgzL9YzHQzvszvt7uHxu1Evmz+H17mrfzMicr8XZ
4EPGa4tyuggh717hJcee1A3Dd+sw8Q/pqP4k9HfcPVEn+pvjABFDG9zVOdfGUo9u
3Phy8W17W4wlsItt4+am9DyksgNbtFHWsFqrUabywQpclB+eULVuC7dMM62OeDqK
G+rrcbPC3XERnS2mGPhXM8be2W/Np06LIrqbBGJahjyJLutNYSi30aYIF5sZGPLp
xerUIJXPns+VzTuUQrMb9a6ILTQntS7MenDO1m8KtiJHkKL83VWbWKKJQoex6naz
MNd0gvEjHHaACcn1wBatuX9NT36/cZP7AVcqF0DmrizfKDk7mXad2Nf4HTGyKfQV
kd8tVuCI4xppXpQ9lYKpfDCiXEzvm/m3K5kwhU3QtRn22WrDZJ05H2Dslo3DX1M8
ctO0OtoeqkXdDLD7BYQX/Q28D3s76Zl3QdLCyViA4P61n50TE69PEN/TWHIyNXiy
yF6kIEqe0PUcAebGgOu2RbvVnxb3ev8xBEXqp7abLJuhJkUVZWqb6sD+eJ5DOGLz
UlUVnXfMkcIOOoN79xh5NTiO8g9tX5WPZASlbNwKZIyXFlH7ZQipEp+3pEvY2v5K
1zlLSOYpSUNkOKjKYCvt7ceTa2GnzRBsYA3eJMQdZD4LKbT9iMJ3yJeURiO/O2gr
l8pUUEmH/otLaHVo3OlSFLVEpJZkzT6P1lP7XoBBMJZ9bnJ5dbo06QqUB7zcerPR
o2sYovzbultRAy9ZmbIdBL3pYfR8lqZTn9cUofHG37vc8SJVY3DEpq68IComWbrX
OjcyMQbTzampkf7TAwGu5NwlxfqFtL2BgMBfOXvF4DuPFFfAm8YhnjeJtTuwIG63
V8rTBVpK9fbzkZJPTM15ZS9Pw4NU3jKW1ENy9sZSZZY+7ZAPwz4ndIgpHakyqFkg
oWt0UxYpMupsaQIdglhkeR8umj2AddZevjErS0Z6X0w2tNNruPm+J2wS5eMvvK6X
J5UK5hOymdUKbTeAGLkEhWgpYwyRpQLMHVkpbpUsNyGwAdqZimvsAWiXwseY2SnO
JGWwkeGr6paJ4ZS0KsEhvUyKW3VFGRoJ4fDYvCcuXXSlYTcH9QGTEZGzvWc6aV63
q43+T89mlZ9xkxHNzDq/LHDiGJ6iJw1CQlubTsq4W0WTwktS7CVIJtv4a07RhCd/
f+UNt1C8hVGENqlh1oZCo6ghhMYjdeXi2cD+2VEA3HqU8AXgPgBqVFwUtPJSyg6a
+xwI+rSImpbw5OLoGGMeiSuxO0f4gfc32KT8i8zQLWK0tJHDdZXP04DkkUxk/x+R
Y+5eKXb8f5bAQd8hoLD6vqBV1d54tC8GDHD+G1Xfslzp5tWUiQhphaaeq5ZGWrU5
UFZWiiCZoMXEOMsPzW2bw35ETKc98KqDMF2v8tFDAKSVdRhPJ/rojwgq4G1v73le
w7/JwXsUdLRMBEWx7B76IDgKXRnDYNS/+8sue4fM4LY7Eefxnm3B7lbv6gDwTYVs
60ZbMpdvTbw2QITuZY0y/Fn358r6WnyENSgb+VklsFmChihakIgilOGkRM+HB4PW
c36fQeM8ELZWLOmU6hk9w7sLzADi5xdD9CsjsAmVwJOkGwr2nQ+zXSaCipdg99xp
/yFncPynBCgIkIQMJ/q5pOdeK4mUPyUkFx+lxeQL0amCinNB/zUTy0uRXKwgKA7I
K48ZYEDGsbigBfJ3cpvygKLzMXgAbkIfJ08BGdNFwcRwycH+4hRozuGgExah1P6x
0xdQpxfn2gAzy/KFM/csLqcHlO1Q6lecx1IYqiKMzVm6sUINdmols9TxTc0Edwjr
Bb39eLOTiEGjz5vOqzLU7qE5I9WrbErKqK+bQj0EfuwvjHtZRYb7NPqoHiLM1S/5
T6aqnehZaRdXFkSJNR6Khst7EL7ccsRcL/imWAL5eSnpXdrLdHdq7GaHjPRxvHFT
FJjOP2HLv0RDnjmzesUy3V/n4bBka0yv4z2myW4C0iLuNZTNkn0Zcxu8wKTePFEu
N7DNr2+5n785kK0/MKh5IJqJvAIQmT3PKV550rjYewatsywngFr8YAXQJS2C68up
qjHLJVjqV8lG7rbpWtVLQBXqTOzAhWpL+Mvp0wtdUG+8ZKiMQMyNlsrTrMLrY1FU
k20e+ePoGPAfmphaNLYQcQ==

`pragma protect end_protected
endmodule



module SB_RAM256x16NW (RDATA, RCLK, RCLKE, RE, RADDR, WCLKN, WCLKE, WE, WADDR, MASK, WDATA);
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Lattice Semiconductor Corporation"
`pragma protect author_info="Lattice Semiconductor Corporation"
`pragma protect encrypt_agent="Radiant encrypt_hdl"
`pragma protect encrypt_agent_info="Radiant encrypt_hdl Version 1.0"

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP15_1"
`pragma protect key_method="rsa"
`pragma protect key_block
Ale6EdOOC/9gkzSbfyRbkGGvlD2JZhvDN+4MgkQmKz1wT8zu0qXRdr9zC5knD1bh
/VmvxucZXSDw4yn9yLDzud496WJ9UMbmdFLqlR5fayCjzy5mMyBdqW4OzLUUEZLV
DbtuEui9f3+o2DW7lq3g59g4fdHirAbzHPpCZy4IJyFVaWjj2iRSimOM9y2LrF93
SVcATu3iBXOMemkcwlJZzZsEgGn44K0TAA7vQAUYnSU0ABkFaSfvWqIGkSMpQrR/
ZBvFK7Zv7RCXCwrL8USEO7gZVfeGODSXnmZT0xrlQK8ElKawj71Sa9N98EImJtHR
71reLGBrF1hPDSvNJyvdUg==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
U62IbQ1fPhE2a1YtmJN9V1eg1g/w/ghPewZGUlSxp7831J9eW7NuRMJ5L+YcTcCb
Mh5pQyUdIHHQA0m7xy4sutqTLz2IfdNNrKvYFE6BsA5ZwhcmgSKMVGOP1h7Z35jc
SY4M8I0r4grwmwYk+EIfkEPlGO9FtD3i6ubfw+wlwgOFRLx34Gqkr36er+4r2ANW
v3OILUCjU7xNrpFNIhm+SlPHcGfoIypDv3+rAhIT4b1DlBOljdCewUMfhZDMBHle
majLflTcmPveNwlhrIk3hQxU+/KxNXA6RmLpoM7grNj2yN/3p8bLcCV/zpRfLrHY
L7ft7TYfwjnap0YJ0gVr/g==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-2"
`pragma protect key_method="rsa"
`pragma protect key_block
J3yj1SD1FVTnVUgjqRtpng/rFTPgXC9PywNHtOV2GLLnieH2n1/23wPNmX0+AIX/
AZRMoB8DYHyO4ywVN0+AkdjoOcMaL8Yajr8hIZiX3Sot6v/czkUTcCUH3Q3e4sMd
Hy3vue6QJxgYqhVIdqTBi3vqegIBe+jCp9auFmZwkppY1FwGLfmzRIkN67AIhbOH
T+ZGkwLIBh1FkoX2K75DbtmYBgu1XpBm8DxEScT3eizhQtrk/IPVG28j+eY2U98U
3yK/jDND4y5G0DzUAqHL6qC4+9fQHTKLeyMVXUsK94TfetjqdZRobjKGg+BPZU+t
UHRtbAXCEivNEdxP0L5kUg==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=128)
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect key_block
0RpozAVunzG+1Zu68lgC3YBlUni+tWnHVsdyEKs1HZhkR33EXYqKE9ssSqAnWx9V
NxVNSFPb7oh/zCW3ReZ2DY4HcSCZAyKbKg1W9UNXMczYNEBtAgTAQqdFrt4eTKut
pbKPDggqTvPmM7i2rOOmFLwxBSGhOYBSi1V2zr1kuEU=

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Aldec"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect key_method="rsa"
`pragma protect key_block
wq8TH3SJsFoHMqCq9XVwADvEd5WptKQQez4Ns1Xm86wz5KiqU9xRgB7NIc3GIrSJ
6t1NIpuo09K6Caxal2M5FMa7MNi19OOr8aZJhD1rpk1wdJl2om5UoOg493KTHXMs
aOptck5wG5EJ9NVzt5PzoIkUaNpOpFYm8K7Wj/Hng3di4s2QSplwkD3gZnf5F5zX
fzfh+MM9SM2upKDYK/VmZQbjE4dUeIXIpGdY6BDqV08T7hK73l8DBC4IGAAVwLvU
2lXooBuM9kTCyZ9wLLbLSuBce/vdzUr0CzaSA9IMO3I0zYB5ks/n4v5P0DX4ngXT
2o/ae7YegF1GS3RRbue5sA==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect key_method="rsa"
`pragma protect key_block
bWC2hnrYFJ+dCqiqBSVY1rnHyeHWe2Qz9IsZuGGb3ZqjL99tcVmlo7LZNHIWGXTx
eZmDFxXt7om/+PtUbac/6+7prh3mNCzqJMcEuZNMbNJeU9XtmHQNbnvcYXqdCSND
CM0eoNEa6m5+M6kwK+65OxvXNLW+sbuWu2zYBGCRVNPEkvBGsuhgu8kbzb2UWSgB
XbhnzUTfZe+cL6vPoXUsHATlUIBfkM6NTEptAJBaWz9ilnxqd8YTWzkYiid0h0z0
CxTnHD0CN1qfkb88vCrLShmJcw/5cjE7j9vB4ZXLCYiHbFtTZrZ3fZxNmNIi9Yue
5Y/JsrlE1Kc3gEqV4kKgtQ==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Lattice Semiconductor"
`pragma protect key_keyname="LSCC_RADIANT_1"
`pragma protect key_method="rsa"
`pragma protect key_block
Q/T2nOQONFfBwdoRQgvHjsWz7BtO0qAHeqwjWrFKeplD7e72goRTByVUrYcaGsCl
iPQnd477AVXt4jOvoRcnFzv9sB6e9V9wNfGQ5IUqgPVmkiYkjuU/chUXOY3ndZW6
N8gZjUUzpoIMNKRp3bqQJgAH26SsLYRWvNxusitm/ExFmTdZNZS4sCHBGeNws/wF
aWAMg7YpmrjWvsDTV8tklUo+VWv8AM7Q4EdlrlCyqQgtXy5ENEl4mGqJn6ZmLkcz
7Zs6/suoVHQ/22t7ecivef1ML3DhXNrnLs+67U4fdaqpxG1gKm1p9AYmWU3fxXXP
0wiOzGaVUDYSch7HFr+X0A==

`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype="base64", line_length=64, bytes=4016)
`pragma protect data_block
TQ+ktI7RFBvvbweXIJp7PjkIbY6uwV32dmhTxYikcFpP64gSfDWDmPU/LaxXgah4
iWD6TMXXzy9ma/93gs74TfeEFPyKGabiLeMq/f+2YfNiIRyULC/TepLyJuMQnWxv
twf1Qv6xee0Uh7cf8ecx1g1FN1OVD0O4cyP8KaNRZ3VOrtMYuh9MIvftsxviGH5T
tXCntBH+Jm5QdxMZWrC3uekfVaeMHn6pgwaLSqr/XAIbFv+boVEhIcAYU0rXj5DL
kKiworvd5lhb+agzH9Us1tD9lU8s7a8vcAnjEFZoMgx4soUsY+wa5gUCCljSJ8G4
JkvJaAOBNV7Foin+QZ//KyVi8rFktgx8cTdSGxleTDElxlvumdZpeZvXjzed8Zco
7t7iPL2cd1ziYYPrQiAYgfdoAPdwBVcqOHWKuPErYUm4ADsMJjMd/SbuXtSbGf4q
UcxNz6haFweTkMSP4418Cbi8Akp2oLb1nrCaFwCllsimCqHV9Gs2l79QjFZoqEn7
tPXM8/qSM56DhWlI11bWKOWyi00n3lT7vbahJdvqn+RLHW8p7WQkjzWKxr/z++ti
DXgNItCtl/57lZn1m887RenGq4uq0ccfJukWnxW2LqUrXhWDrh2kcgiurVbz6i3H
7fH2wh4O2URQ9C5oZrKzaOGeyzZt3mf3E1jb/VuDjNs22hYZhwV846V8RMJYI5ft
f870kgI/BlkBad5brLMQgA7XIKZkjQkVZEfcXbekvtMI+/KbOqp+hnjH0AY7GBf6
V2eJfDcEF105VWnnthMRQJrWSIW4X7FyDGaWSS4/Ms5a7nGPVfU4PtrJMzL/LNhO
5Ic4x9Afg2qZx26mLspTSqNaLnoYzPOS/SuUFx6TNV5APoF9GAfk46WxlBfJedQV
2Dh9FNuMiT4TZAwifcTwPxr0oeKAfnAm0KaYVdMZ6SqjLdk/8IhII+yHN4I9Vy5Q
nSpGr2vHRaixPCIbizW53kne3groneoh7Jq5zmfxeM+nrNb2ggXgFOy85/SEUkmt
EPc0twqbop9nremo13K58vp5ku/+u3DDor4yK7eK6zHCDmm662alyhmZj9e3UwpO
eiNyoJrse2arNNx62fyIQwob2XWkvaRcAVNngWqBOLDrWqnR6zK6J8PwRXZ09LdU
urwAoB6WVVXN0BDyGWdGttUTavhz2dOejcZm6V9nyOZlNeLzf+25rS4xBpBFe+Z0
y8u84tk5gOL+KxCnHR7mzEbqhNPXj1FFZITXBmgD/asKf1cOPPp/ZSj/IK1P2Hmt
ydv1bCI/ySnBL0ahuucNipHSu11younWrnZAkT6yBtreEY+rxlxuOA7iSyHlaUdb
VLccwbBpF7zISaW1pNH5kyK/9C6ZBFa28twpXL+RlLemyIc68PYndYli2A+lyhRX
DgSzmKayZuL2m0zjdwuNLiVKSG7mM6fBMDq5Y1/ktjCkKF2ip+KLCJsTVPYxpnNd
o48Vm1x0c03BlBxqI4TgWcCzRGJr1DGd7ZCDrEfmczTwNksOQYPTicdOC4a4N84b
L7kmNdblwjFRyqS4FH7Yq4dEywnak4NvpKp0MuBBdZwn1cRjB1DOzgNr6CSuW96Y
Rikh8jxzF5dhDmwQH4aCbhnMh16LFQtKOfGwR5Ny/KgsCbYwsqkueMWeW0+qMgjc
Tqgqob/7QERnUq3XmrYvN8YptrA+9gFlnaRpg0vn1ohe+fSCzXtQcFNAQzztuNrx
sOhfcaGsm1MmLiWHQ4FGcmsshG0GBd2WOwSnqrLBWfRpcHxoEK0Mf5XIaQXkCgVU
USOgqNol0RRy8MO1j7J8HfZNPBoZSgnlwVccBomzox8yST27jSjCxOk2xggA09E5
jdIQYVL1Y6FpjdX91UDPBcbSEotWTWz41+WRIHGp/yMa4DZo3PYE0+e5MKKtxk6k
oVE4XcNn0toTY2MUaRHUbvrHg5qbqDpcNQJh2PuBSyCZjpTxBy+P34XD0d3WTrdM
KpCrpfVmcs4GoiF4rGaIpuNujNeyJ633dySU1Q4C6whsWgmMsFinIJjR3hN0071v
UPh/FRnSFf4l1OC1K0mXVTUm94fbAuERcRPaJOs3l4M7SHR1QvtNv5KvKOYpjX9k
kfW7I+Li0yLPGZ6NFJvaC5zS7DGpfMxl/Ld8BoVRuTHVaRRa9J1H9Ksv7GgxoBfB
4wW5wXDrKB0qTiCh+X58huEkUHVIOU2PBC8lF7XXbb3ErbvbSUTr5VlFh8z6NHz8
5m6i0LRy5PQk1st4Mp7hPLnIpmkp8jsK19BnjbfebXXKBlQUJU1Fm0oo37XrosGy
iqZPdPUUr3VsdjJZ/sCfgmCDJhhpWCG1WaOYFjDYjbj0JGqXkQ8bVdkkwArMfGDC
cSXxdtsZtgOOAdOXzSvBcMaIuZTXXrhIdEqpuVHQwNDnBJsUWbF3xqbAD2VITkT7
gO6Fo55rHqC3xppGvPXljJX8sfbbrIlexxC2uwIIog2lT3sgS79/33AxYZcZ7Ka6
Nvlbe+24x9chmcDJw1kvYkGvTQULSxsDGg1QH2Y0iUK2YXX6grJSiXbeBJn2sKhS
0FVYqJcFALNKzYqsiQJmb1YyY8axENuvrazUPMz/jQRA8wbQ61VxLY4abTnE/3Ed
IJrvXBIweBjoDt5Wlk7uRWFlr3BkrG4gWswqhAUNu6isRAHTZhWjwlJuQ6rFtYqu
nLkFJ3PRU7FqLdMvVbWdA4uE8+FQKK84IDTAC8AT8lNl3+bxvjFJXgjlffrrXST6
9hVkv2pUZZFMD2FNgo1L2R3ad79pVVWPRDb65Ah86LhAHrGFTt7gPfkcXoEZyPPP
vmoo3GAwjNg47X4961yFSNQKKHbusiTzKRxicEnYA5bKBzboCpKUmKfggMo/SLnL
9ndCmq4f/+tlzrcKv24nFIV6VlR7oRqERA7Nssz9d1Mh4hltAcw8wCf/eoT8WpcS
a+tdwE3U/woaEXmhJf9As9xqyat/NHudU8f2g2cfq2fwH9tQyPBroMxSnAtE7TFV
8a3DOkC/yG2LtaPgvUXZMgeGAvdT1HjjHjekRWuuCwk2QrUFD2c0KdnM4O+b5r49
X60k5kG+6eBEs6oz1SuQTsvDGbw76to22ifDaJ/kXmNOdKQxXh2745XJcxtesPAK
adWIutg11x20pdoMO/OCXcTAHU60QdVOokenJ7frHV9jt9Qcr+YlxMCrHjkK156V
rpP/kLIImKbYUQmmWbFtdKsVlJXRAPpTSzYNYqkh55A7YUndQdfizhGAPvD4cT6W
NgxVFE8PtpBZGut121rd6TJtqoSvZv5P+8GG2gDI9I+gdrFhObUGE0B7X0uUxuv1
qhdt9qyQ6qpdexpI1N68z62K0vVW+/tVc0gaG0rrK+ASbk1l4CJwyXTg2Elxckqo
GLw7iX1sB4qhJVX2qbQdOTEyo1rvTBh91EBLKQGKRxSn02okPCad9nsKZuxodMzH
CgRbl18Kk5f16FBlSzcaYFSyrIrisPd+f5bZfIXFeFxmNovBxF6Jmh637KUyIOM/
204ZzBzU9reK1gsL7yAer2waklDew/urHPY+30LVwwIu/tuGTfcw8Sw/k++x0d+n
KaaOb/LK2mT9YP8bBxzmHa92N1YXLvscKHfXPCz3mNsmRPW2rY2P1qBKYWtHr/uh
VAzieLVEfS/QRghVFu+ZUlTz4w6sqrJKG5z9VUO6JzyLkKZdx81/7yDg1CL7R5Pu
3vGiavXFT6SqEN+TBJ5weRYNNJ/3Eh2eEeQDWFFSJC8RZZhlT8vYvWvsb1PvyNRC
4bZZrqC8jirbztUN7BDDqRPzjaw6JbwLROezmqdjgRp+GfD3V58DmCVPld4Ru4dH
OZQPvdXHEu1vb2LcbHLg53kgbmPpKWlX1ExdgyygnQSZW/N9/aM3vO2qu6rMfs3t
BUJBtD4tvicXn+qVSxPFwpheH8W9uUotFWD8BfRtmhS7bK8KXbVjTokVw2cTahBU
XQJ2QLV2XCjeUN13a8YsOBKQ13Jvscf8WW3T5uohYTrMLuIdX9AG0W9J8PZnpm0m
V5jx7V/lmHaG2wwouDDodLQNifN1b04db/w1SklFH8YZlgDv+PzmFwnehC26OWhS
xK+c8d35awq3gB/6CrDJod2Lp5mBy4z54sc44Cgl3MJbODDQ+s4DtT/VflZv2YAA
QM3G1tPQNKQlcnv5L+yJmMVG3qot0XwGlFxueKp3xZhEX1L1oKoUAqIHXhevtk6t
cci6RNnBVT2GTjvup0y1pRtn4jLaGPWvNjMKlmPdVWNRn7kjUpYUQceSCFMGRPJx
h4EPW63AC9npZtDHb5gLGf3Z31mRmw32m6dvLxZh9upI9RCboMDmjWicLX50JXnv
jfMqIXS7dJiXlaRn7n4g1ZMZzse2wY2f7yXKlBIdVNWbVBZ05m3hZqoKL7PXU+Qp
BqGux+5zO+d9iH9NcIUlhY5A6yBZJvBX1F4gMQOadUi8Wxl0rBuJo5HITvXTIy4b
rXucgoO8t9n/FQR/nsMNzNp23VECTVqGuA5MDz/+R508zmSXcBQfjns3m5EltxZ8
9oxqlCOEIA4gJNwJ3d98TLhIkjFvUXHgkUyHoJ/KX8DdxOkqVNwEBwAEswgsC+r7
AzGHFpfpAvhcKlq50yyXXNUPm2RBSlTeWLLKo3f8axKAZzdZo1bWtxgbt7kRd4PG
nsaE/GNzfgviKkOwdviFWa5qlTxV8sRSp23k6DHQ8GLi9+nAC8M1yFOrUEjPy1vX
8bMwQDTfqZY6OPw/9e1p0BQzTxGIVxIuKOUMeMYcBNnWARVBENqv2J9XYlo1TQLN
Sh/KIUjf1AVcFtQq6auI7cqgFqtLVBlAIZJsbEKzPk4548pmYtODwZbpLZEJAePj
UTcWEbfAtHtlTU2pYPCY0W+r1AgetelQxTNsdU/4sbW+sQnMnmxkxzmStP+tr4hN
1R7KaX1k+jpa71zH3aCEG1CNnMq18hNLKpvcpHcyrC/x/Grhhtd4j7zMCh1OHu4l
8fapZEXF04xIFTGHuQf4g2mMCQOzNFWNpboZsVB/n+cgTDRG5S5/WlHGM/5UNwDt
r0wPBpJZnQA11Ipg53cER+s2nzo/Hcjp3OeUPTkJhl4n7i/PvqmkB7sBVT/c3C4g
PxMbhgRRSurSA+bzxdLZTNQMeiR70VGRoAwuHODfsmdwFGzvcwEI1sZswv89b+7W
O22wMxFl2xDHHVgLNgD34OFMU2L6o0avLVLQVidhVjYSR1N7ZYd3EKnmgkc2IpnJ
pTIpXV0lliiWPVwHZWi02UZjg+iVy1Ou/vGAUn5pBYGRa6ibDtYa+Uj9pOGbAaNq
WbO42RdRcKYK0q1FYVz780j8Whpj4/LreXVVKcff23Y=

`pragma protect end_protected
endmodule



module SB_RAM256x16 (RDATA, RCLK, RCLKE, RE, RADDR, WCLK, WCLKE, WE, WADDR, MASK, WDATA);
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Lattice Semiconductor Corporation"
`pragma protect author_info="Lattice Semiconductor Corporation"
`pragma protect encrypt_agent="Radiant encrypt_hdl"
`pragma protect encrypt_agent_info="Radiant encrypt_hdl Version 1.0"

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP15_1"
`pragma protect key_method="rsa"
`pragma protect key_block
6vL2ajSKwGkG8F6JJqOERVnft6QbmLB99jnFsN+fwwaQC5JYJgv6yF8iDfgfiWeZ
jEcs4caGtAfX64Qii5h4YlnEYMsEcfQeivzRStkB4nQ42iroaUe4ZeFFenVJcMV2
pBK6SysRrzRyeDOdSo0TlQCry+m6jJHNbfyNcKrnh5d27ntF6wd/FYiIVVEWfy1X
gxxqyylOa4XKVW42fcV03s54KH6a/lZctGNHroGa1psQubXqwQJDwdS59l8B96Ph
fH7OWIJJWW26XHSIiCF/vW3ovflOnwRFqw0U3lfuT0GCTBIquBpB/M2259ztGAPD
jhbP9lj+0noD1vMe/cQadA==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
E/79d1C3DGJ7vI3xSISEjBiG6yr1JpeydS43d0FmAgzwbXpvAR/71EsgDB62FlGh
reno3auIElpTLHxWdQ8FGn4mbPUaVsoymHOzTrAtPsuLGsH6SHUIjdq9vfkEuPoq
ZajxkBOVgX1wzYd3nMlAFBweKhWFznX11jr+0QJOxf2gl4URWE0mpCU/NiWocMSk
XY9fBn5p7k2HZr3WcG26oYHESLGKpv6wgmuVd9MrvLDjgMzGGIV7gJzq/ahcq5uj
ERZeVRHZKLuj0WNYDlESMAgsiagrXq/1ISR6Dcj5FlsxD3tMUnyrWxX5kc9XP9uA
syHd6c+IkLexpDAzuhlJbw==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-2"
`pragma protect key_method="rsa"
`pragma protect key_block
ObzT4SId3IsxGIUouZyOXQFRh9D7TrYJEoSQbLpFk7kInCxKFOa1yHr6HmFfh/BO
pMtLbcpzXAUXI15VbIW/QJxf229kg7a6r3FY2zh14y2072UyubRroRkOtbRHo16Z
407H4DcrakSe7C+jToGaF+VWr9SsHofXn47U7tDU/bI8nF9OUIAvw7FZy2P0Yogc
TZ48CRd3hRMTZQpTyBmYyVmS9yd2vtlpYu5WFMrTSazP7HMM/TjsD191P7mc+vMt
YvAbIh6QGAKSToQKB4j34kiVtyWsVp5KAc1SNbvliYsuMmuFBaS/fYQmrFmwfOUt
i/1ccz4Y/tpipKs9jbVN5g==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=128)
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect key_block
ZhbiPRJpZjuU3LIG8UDyjz2JxxRjBok17MvDtu4Uau65uIB92j15bKXkpdZhffCs
FnFegE/x+cUEbIUih2Hk3xw0s43Lp1c97viJ8+iL1QaopyUszO22C3WeB3XvRpLS
WeeKER7gGfQ92SGpvVN6hmCnrlV66wcn4boPYxOkvVY=

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Aldec"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect key_method="rsa"
`pragma protect key_block
zCGB0cIeTRJ+0eHpiOJEoQj9Pw1Qcbo/w5ZaTjA8qSI+RWA4hepFtx1iIUrFbG2C
puMercbqfWOU+an9alqsrkXWz5lE8ryDwelBwKo6ZElyiIBkjB+/HchuxTbRlIZ0
f7EtugcEgPu0yoLdLa50k676NCMKTlJ2+yPm6BRI1zScTKd/fPSjGooryXAKjfn2
E5+Fk77Jv0S7PC9scv+e1Ivb2Eahp6Kce7sDISzrHxw+YdN8Ed7JcqgeZA1l4tR6
MPRyIB62Ec7H9pGGh5gLw37S5QBamE2YsDNmNEf36/VcdAPB6e8a8zB+e/sxFRpm
yBbL3KkaMMpihzvGIHT/Xw==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect key_method="rsa"
`pragma protect key_block
hCDBmJGmqyGHPYCsP0T/dPz+S4SiiK6GThV2JN8NEWaoeY6MQhgm4PMH5My7Gi6Y
/b5Aml7FUvHOEc0K2pdl/8MzZzXFqiOnL9COkpd12yKqo11Xj9r/XRaflRimJV+Y
aWAl1x1VDDUUZdgEzUIQlNfszJSXnlEKx9Wpd64DX7VU5DLvosR2zAz9VJcrtJK7
VJCnHyUEr9fN2zWm2KPgxWOnkEqzt9kJzAAO91NG3IP2pq+FXqb6u5GgJmjO4z18
I0OUvcAIbEyj3FO6sX8YfFKgRxrkW/NujpPgwKjTz/wE7lKJgthe10E4ns7EA+Hp
2dXsTMzhhBpdtZmCfHmzpw==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Lattice Semiconductor"
`pragma protect key_keyname="LSCC_RADIANT_1"
`pragma protect key_method="rsa"
`pragma protect key_block
w9jJdsMjxOAHRJ7O88rwu8HISPFrpCPkuEIEUgEc2TmKYqUBxY7chGvOuQ9iXpYL
gjQ6KbJYIOJ8ltGATffPgUCW2RlTn3ao39bxrDW6xfZcCZN/QrZr+j19+HH3oO9m
T8mc+Y3KEguYtNArrGYsz3WiL1QZsR41+2pTy8aG2UcZha5o7U0qG0ujn24RSc4I
gKbHM5JQ3Ux8JCLtc+xEUX6ZsTcpd3SXxIckZrNssHqIPlhwxcbxvnHD4FvOjOdX
IfF/n3RMr3nSFpUH7WErvjnnlEQeN2+7LlRter1C211p5Kv4vVhw7Ascx2bV/lpO
Ed2u7pqdtexOlNWRbOupbg==

`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype="base64", line_length=64, bytes=3968)
`pragma protect data_block
01uSlhUZ8UQSTHRKcHXh1WxI4efyVw1rOtPstr9EyQ7BdVPFAXY/6qDFklfXvWRo
+Dy1wAZqhNRX1tKdKomgRhL7R00wdNJE1ydZV6KtDk1UBw224tQxIZZQNTWshQW5
fk1KINnluf+4JJpLG0Azb7zsQlk8BcJbN0HK4uqI4b5oMD1N3pyKKy5kaO7n6MsL
bw8OXSDG1YhQWZGIEAyHEvnP11QPjqFGAIzuPv0SbxinVoLU2YTuJJQ0ZDUPSqEu
TPJ8WpnQ+ywjqgdklksRKngFgAEcTOmJvdNETv6FbaTHdOdfeTlUxqbve4vLV9v1
UGN1Ym41GolhpUeLZlbXU+EjA2cAPJheqF2UZD+STwQM1GzWe7Lxd426HLw8Xhky
ghAm6xZPQQBavdO9RvYyvkdi8j36PSYNK9OIrbz67JgWffl/UgAyk0zM93CWFe1/
uB/mC8IVP6aIgq7sYNb3SB/2V74xYIYQCH/4D5YCHbn/VinemPNNrIG/aYcn3+ao
U49Zqsh4HmmXH/22WmNKIu1lNRPkmaKg1NGG1AP4kqKYXrJhWsKC0vXOiHc1voRl
b+/iFu+H22kE13SCy9z/KXLyZ9vKUsvvAM/oInkUjeigcX62LqUksHmJDjlXTHE0
uouhLiuffvWDVxbW+B9179MrH2Kaerd0fWwOM8GdjfqwwTITFATJlhltPCXvpDzJ
OKs6GsVvHtIejdv/vbQsPjqXe8admwsOrJPzrch+sHzFhPd4N8K5UM7mwYyaK/RO
JRpRKC0YatkhYLgL3VU0fBcxMONrFcFtQ2nWjr4HXg1DqSpmU9VTWCSpHLIhd2gI
NONHBtu5UdyMfjFoJrirW1GFFq0RyxTxiIIBd3UtAZpGjmJ9Xbgb79B6Aqm8mPNZ
z69YuaGev4MlgB+Jn64rxCUvA7HUZ0gEozadR/g1ZgKuhigAJ60ftkGm5QAKoUBC
KsLASuxCgvK4Ukq6QKSsgPuKfW2NS0Bj3+KqK9sAMtKyDb59n/a8MprsDUo11xFz
ReHAbLd5Lpzer92FzxOKoGdrj7Ryvk1OJP1W+deISUlQdcr27DIAtymJDT2CGkTg
sdmdQdeGb4M9XSFha15N+uAg3XPYS5RUyaddDsrZ15ixvZuhxFrdcgAvYwptiN4+
ZEg2QrWi/NQTnU9N04GQkLZyYSsv7LWWqm2hGPq8RBL/tiGLekk4wlxOf98AhXPH
yDhS11SIq1AX+FtjCxahr+PaZlYem9e9CSEkX27Xc5hFr4qblkQo0LGOohxRS8nn
/zBxlWKk3xoCvn4RyAa5baS4luQXFdUF9zlISI1BIfw22Bl2lDDInMwV+3Cb65vD
pBBsIw5dEC9UFn9zlGERF5iUXJUGgFFmCF/Y9R8ejg3wKdpq4DcDpdo4j7rT1pEk
4Kl75lCcMTYs7JuFBgXM42Jd2v9Pdzw64qjVrQ2ht9HEkT1AwGgaJBMoUq2MhQlg
xs46AmJGSoKZ3TUUqvZu+4EbhJcnrDIkAs3xH5Z/5KczeRwMDTSLLic5IJcdLEuV
u/Nm8KHxe7rk81RkA5XhhLALGYYDPlI4YJ0w1eFj1vJMI4KSMmVnXRPwoNAwcNQD
YSPvXc31J8IPAMTTw6qKUoi0AzrPvIgY8IdJ+2Z7OpJO2dy/S/onLmpW4DKUpHkC
NbrvH8UwZzwPE+wQssNH2N4fjxBlKdGYu6HPq+HA34gOugae+ND2KQA9CIhaDdsG
a468Y2LwVPJ3UpsPDfVOLQ9NlYoYVF/Dzjt1+wBrpV5O6a5ailf2I1vyCG/vUbwS
oR9VWXFDe72rF366PikbW0Nz8SpjcMla3ME4ctMaCoMjQqVq0xB/G4Qm3Ux3Gx2C
RMrNJyjkgiMQcC2tpztAdnHzBVF/81Qvx1JtHua8zrZ5WwSuJ/3iqIMQv9bbUuLq
i9N4KCIm9fecjlA4tSWWbFuX3QBc89ur95Lh0CjULfZaJGdbK+//M0am5axl8CIF
HxdHu0wa7miDY2NzAGB/YM8C2gv87KCa9STQObIaN9yFr4LdxfMIUZAJSVWBHkmR
OKpaIalBwSFaepePrZohDnvQg9wNneKhxgEzAgWDoSvMNuqfGYOt57JA0gvjS88Q
G8gpEyqMaBDYOhV5eZaYG8wxB02rSNqAZjDDbHuoBknyU51qsEAZyOaT98aIw9GC
XHES+TRCjZkj84A74emLU4fCAAkJm8dggd760ryzqIVpxcbzL8awUc7RWRJvCg7j
zD4RXy2+CoyV36B/pvs6a+IpxWvOt6wtv32xQ8sxullEdbROEVLId5E3SnQlIDff
pQhC02a5TMtiHX7J8XlfkaYKSjTKsZZ3S1ylfIueQ+GgTaSZs8euIzinr+bHxbeH
Qu/vaPFLnGyhEMthfzMlhco3dKp3Yn/Vz2fLwIer557bWdPl8bYrr2wp5yMZkIdT
2Co4QvrDq4YSc+Mq2Ex3742j0SDWjB2jWuFh8bAkO1XO8u5r4EIxwV0Rv5IkZR2o
i+9+0EBX/10T8T8IOlP5PoLxSyOooO1gYMUiEWDdPN1ZvggqR1sgSfenQwgWrXq5
i4T723k0akgDqBFhfQGQHgxWk5274RapTYstQNduiPZvYxpskHwCnUvQR1qI7259
A1GLDJIl46zrTSAEiCpqzFfIkuN0n7PY+DafmqmDqpy2vnv3N5kfY2exRAu1fsgk
XnxjQkfCNiI6KbYLeoMZ6jgS6irpmOxrLwGXvAyKMGRtAZwW5vu+sm152mgTFcuU
FqynxiqTKrA1w7Uo23vj2rFywtF5TotiWjSselG7pVoG1Dj8a6F6KIJbR52qE7p/
MQ5MFlaa8emBIs8ernCxDcR7gbRQFz65AHNo92W4xoF+X3DxAME4l/iHecqBJiu0
+jPvZgF/j1DkjFJGk0z8MeM+/KeE9gimUofeJvpQsWOC2ijnddQ5YOwOyep8qUHk
Z0uoHuMPUqoEJ8+lq3uY2635Hj4lbcTmQkS7kGP+o8p2Pl7mFlwO1XoWClsS1IK4
kU7F9wn1whJq6BKGsjn27msItnX7kZsVyfr2zvxjED3jku6By8Y7ICqgqwYP0miK
J+V4t40izYDdzhilAM8oqIjdMBakWzCbzc1oTDqS1jHx/WSuyANtFiKYX5z1NAIe
VlBjyGtZ7qmwt56tBYHp5pGAKVByPRPM+uUKERxWKRUTe9hkRtCb9jAyeEbDyxac
m2TCMNAbtEUEEhXPN6EM6TQw/HtSd4b4CvWoSy/rN96o/BQuvWa+M4tbMdqr0451
vjZq0l6oDWUGBdtQK98JBzxs9PFl57iEHukLL/LxtB0TtznmT/xmCzW2Pi2nhq1M
FuP9wxjrdI2714zp+mAY58aPEMt5C8SXZX1yNrv0Gr7MSGA9k9cohkcDlTznV5OU
MQL/+8kxB1m+nhtdYn+yaaSwvyG3tf56IjRgB6DxS8kvgbkvKPCCWmr5PoYIedst
hGoqSQv/3ZcaI31LBDHHlBp0C3o3w1TCRog6+ZiWe+C5Xadns4Fp/0B/kr2hfHKn
2CUHfzDmAqezNBCHQZZlCY8chqeMi/3y/jXCa0j18KlWRhLHm52Cl4xz2vqVioka
bC1s9Mvds3C12aeHBTejF+PFGzYky3LuAK8OX37SDIy3RY5TLrKu0jrUbHKWgjO8
/Dwn3QTNxZheGvCVTc0NM5ZLRDEfvGhTpVRAfnWedb5O1k42zdSAU3mRKJwE8pek
/8iKbFxHoAB2xw8KEdWyWuwr5Auh3o+qRQmOm1znfmHqJIiAhBgM4FaUitpeo+E3
Qg7y67UA+ovK5IrVt/kjRVySotpLMhHOn1u5KxiotmtYQ1T1JYT4lXcomXDaadAy
jHMdWK4xnWZ2Yw4cOmEJzaauZc98wJvC5xot2OBzm1mdO5nbolqbtPqa2LsR0m7Y
CXAmzeM+RpPi5MjEtErDRe2p6BU/mfqErHLsyskyXaNAk8kDcxSVkZlbM8slp1uH
mNBy0mGGxaV4CZHed5o7ykhlMcKalQLjeXgRI6c5UWj7ITrpGZNf1MslOgS2k56i
+VPUV7JzRuw4KQQiRsXw1ba60wb2yFEwQdmJ0Ys9GXT0Tnb/O11jNwXtY2aX0JzO
58pm4a55ygj09tCBa15DqWw3uWsZsn6hG+qjCqnvmLTF/9loDQSn0cDyyS1ZBrzp
iO0uu6A3FB+FAV2K2efHKN4yWJjZ1fPxGtuvy1Wqe2nI2YMtNZKv3VoVKydHsn3C
F+9xvF9cbSnq3AnInotJPvcsX/rAeZ8QM5ipG5fpMCWCkumv2m933EvwiMVMJvo8
tPKbIO1MFpBwbPXhm9TN3ceYDNwC61p+a5ypsTNk7TLE+bJq4gsBa+Ew0oJGXjSi
yyVRGBYaCq1KQqWhnWNTovqNQ3QmUdlJVWCvbtdRexNelIltbhljOJAvtX9YPKdu
C4YyPRchSZTSJQX572B0aBxeXZ50+GabMTjo9zkKBa2A/aBaAiZFo7HG4myn1Cv9
AHiKKd7upsqKhI7gZgtmK8/fS7v9K2ZNzqviPv0H8ZD6A1emuAwY7hDtvw6DQlsJ
7BHLE/sLGLWVyDOYHD7R8+jesWqV8vimZ5Yo91xrwxHw2MEcaazpnzTzzO5aqaWH
wffOfq7yy7aR7S3C33Ioqr9f0PKr9ObduJF0KJeCtnEG1NwRTjDBG1fgklYqp8m9
cPFYd29rJNNLcq7PnhoBJjZv+znV3vwRrnP05wGuqbqc4aUwkedpn5Vz/G7S9oZU
f0BZ0/Jf1T/vMjRPd3ZMv8J3rL/+Ak+Ya2r0aaz6PPm0PJU3zEda1mW5/OhF+IQ8
lgiuXF4wN1sSv3Y6gJWo4pb1yH8FlEkcxDGM07gGEjITE5sR3XOzBtu68w+Q6hQj
I6f7Ty4IfuB3V1d4f0FqZa/kQVf6BFFYuYi+m/BFeR4qioaBY1GuMQ/bnsJreD1d
ibsT7KjWBoF2g6Jv3NzuW45fVujgOF5LikrlE4uK9m4u3iYaXpwyZMpvfWxx2j6Q
y7TUbzRjTR7i+ulMlSSHadOQG9GDi6L1jH6T9soX9DaZ9bRNvhykMienG/wSRkRZ
gGbHYW/D0Y1Fx7AffKz2UiX2NzzXOITWRn0Dq5O4rSSFO84vQ1iTwfTRiqBRz8/C
Ytb3ghW4bdktqlqg5a4uHI7426qLMH2sNmDWkM1NhrSAuF5VRtLZ8nHdzPu4iLl8
HWx0iR+9L3N6VjWZ8eByGsQ5K6tkTnvY6Y8zy0GQr3BabpII+BH3eSK0wyzs8rxO
HUWV+sY2AGTdTj9ilSEXg/e6lMyVawaZaOsz/2PnjYY=

`pragma protect end_protected
endmodule



module SB_RAM512x8NRNW (RDATA, RCLKN, RCLKE, RE, RADDR, WCLKN, WCLKE, WE, WADDR, WDATA);
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Lattice Semiconductor Corporation"
`pragma protect author_info="Lattice Semiconductor Corporation"
`pragma protect encrypt_agent="Radiant encrypt_hdl"
`pragma protect encrypt_agent_info="Radiant encrypt_hdl Version 1.0"

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP15_1"
`pragma protect key_method="rsa"
`pragma protect key_block
JtuevK+zZI5IZ0an5Y4ONHbA7uH2/EOVfHGuYRtb5VxG6no0AI+4Tb4wm3yQYolK
/QqUbAtWbeDsYj7ZlS26fNVoCKIScOzZpyegTrfxS0RmNqjA2NIjIbQq3R6y1VOB
XVHl/KBsORV8w0bd6NNQqsB+Tlti8y/AVrjXt2aFKpPoLL0nDJXejgjfPOQ8a13h
+y4OIzf3Ixqi1ldZ2+gvw7xSvnJHY42nCRYz2d5Mv4BYQP1OM4zANJlPJiBnazCg
SUnxTLI+qgay6OnOH/3pghUjjCft7q1rskUX2XcQqzDGhLItCFzV3WY73x+BISU9
fFx44F8BmvSFdohp0jp+VA==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
IvKkA78bZBfm+lbhXgn9FX+qIyyt+KSR9SddUVDdkf/XiL6rj9gSnTzVO+q4Dqz1
oxQ0OMYm4cdyaYasTYdUA/lsRm5r5iyGbNvBZwCeDExaNm88inNwVhyWMY+F5IaD
YN+Lj6yAuv5fv6y1ej2ZGXd/beLPpuy6v03RVaw7heJKSfNYpJJnzcm62SX/a5VQ
vJa8IoSawoTb8kFa6AC2gYomoUtzP0Rurqaodco5UwquLAV5qBzuIGSq4SaJCQzQ
Un+B6kzk2RLFYfMeWlZ7lyi8TE7pexLy/jnbNTAimiFmkZWWs1uoQgeHZ+saOpV1
dNb6ixFQloqKliKfBfyGUw==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-2"
`pragma protect key_method="rsa"
`pragma protect key_block
fVSWX0iELM8Au9qBuo96Ha0reSe1g0oN08yjTm/rVT7L2A+wVXCbhrxW3y8/ok1S
A0m6f2PD9Jj5oyIaKulnlMVyXzp/AXRJW+719yMaTQ61LugsKASZyTAKw1C40o7U
JcL7p/sxgs4r5hUPSAeRyR9QudtCTkNQhWEUUhpjBx34846vE2JATZa+DnVKrhr9
vlvhKGSFTxOUMSnUFuXg/sZEmdqD5DiBZZYGKZbEk6RRKGL4qZ+4Kl1eNCSMkYwF
ksoI3LOx73nZ7XcSGv1kfU4vnR8ab7BERjSttm88QUs0BKFeQ1z/tf82xPhIh40r
GyWsOLpTLCqEQ0pb7q4kBA==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=128)
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect key_block
BGXX9jjlpwUQZ+/rDQaqLnwGzx1uH/VaslfkgYrcLmRgCohLZenZlEtNLcWaxxe4
M3ZadbuA7ikq896y8mZZT6b786jEyS072XlVqJSD+ckiWMtCLAXBf4Uzt4pJ6rSa
+/Tj8TndwLd0yEqu5gF7rxl9N1VhrbInmS4otqStcuU=

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Aldec"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect key_method="rsa"
`pragma protect key_block
yNqVF2utJoLQvFcmK2qSEyRoz1h/408QXjD0Z5O4VqkxYx4nMdEsH9Rjsv3Zg9g1
aSxKhCCFEKLQFlyTCS/WDpZ0rG9uxvJuX544+tHfJuSDsbkLAlq7hwxTUdfTMGey
fLuFIuMGqXrIje2ppfRZnQOSApGUkcY/YRFNPPm+a1gGKOl9HsyoW2XyebKFPrPw
K/zNfBNY5xwH36jmzHscj4yfbKwlQrOQmNfIUUTCBgHTAfzSXfQ+NfN55rJPd+Pn
ALLpLtGk9tvUcMcNlI+iQEm3UED54YlSjicicMP92hOlvtP1LFkLI1QpCLhuF9Rg
Xq3YNlZUFCSu58D0oJ7ukQ==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect key_method="rsa"
`pragma protect key_block
ZO7aTD1XuYE9/16feQPA+3tyOUNIXP8/+XutOq3IKgC4c7mz3Uk33OaoZsPTgJ9y
XOTMT4mZHW5E6Yx9yvQeQfs3mMcY03x6bEquhD1h73rYr63pSU8yFisW5G1a0+Bf
PUxak0WSnvD3rYMaPuVt0Eb5LJFoDi3JOojKjdBRNHErd/dQ+KTEVf9SFaHc4prD
tbZOYcKNwM5iogE8AMmZ5ZiDSaAS2/B9RzuUn4D/QwU2kDTPl46+FH7JXa7rD+gg
DD2h85LmVUqFUBMsGGVj4TuG/WiUGLyZWnBA6f3LzmA09Py7oBSOD62VbjqmA/Z4
DP9EHWfyOj9heRC1KPwo4g==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Lattice Semiconductor"
`pragma protect key_keyname="LSCC_RADIANT_1"
`pragma protect key_method="rsa"
`pragma protect key_block
YcYjIjhXb5HU8JrqlM1RVL+LkFPj4Xz9iuYiCH8JkcQ9Jy/Xz6NPgOhKDxXVF94Z
MPAM09KQz1O77ewJJPt8UVt4BqBn9tNofY37A2RrDHqRshM8YhG6lT/Kde8eumPG
XPG1CcYtxokjW8O5GoPvcHUqVJy18vJ9EY103abCEtvfgSkUs9oAb8AR+evFtQA2
9NMXOwkFrCkgz+s36h+Owaj9Kzrq0GNxehkNzOfpgvACxXUF8cwwGqyf8q6NK0VT
5YwbrttaO0/Bv3LPVltroM9PVQs9ixh+RWT82kTQGsR85IDAWSfJYKleQe5w6pTv
P1J6ZMtzWQ3X2c+HVuH1qg==

`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype="base64", line_length=64, bytes=4048)
`pragma protect data_block
zQ54vgIuGEFXpk25XEEq7/3hhHHjK+UfrdriTm12ht99L1dzWkLu5/UxVs9w8A/I
7Vc5zWUeY4T1E5pb87Mw385/AGxs614ZmgujYxJy1sRidZApquRubr7j2Wes4U92
OANr8NSF8Ih72mnt1IKX7VEMhKImvJU7zJoePcaKdCXEq9KlHK8fI5BLvlk8QGF+
7vUmJvRuca30ZaNHv2eMDQHtopP3HW0oj+j54DOWP4MFGT0iObKSr8qW0o5sR/8W
DYsWFRpoJqx7ib5usCfe8VZDT21jYSJdagsHwlvd/CCZTY+lxH+qdyU+2qOi1OC/
TmdRkhvpNvFfmtppfc9V4w2nhBAx4+tHKV5bH6XEB7BMqfqzq/rjUBXlQDUNySI3
IiaWmm8YZKooUWr4Q4JMS4JBmSejjwTgynXfQpihm1R4BPq/tvAFCeGS/2DDpMVr
Tprvr9rqN6pZyT9fxiZKeyFN2yVozrXXRp6NrQJjf/ZSNJ6MNHhJvnD9H1D1HHqo
4JW86+TjEZHpIFg2elj2c//dIMhUAiTGpR2KoYveYPLj6Ps2hXdY4XHVSyy+x82L
c8VBj9clUcUkw0lrKTGxtY9qxr1Uq2q92xir/+pQowYhhs2ZnExBA1iMEn6DD2hQ
VlMwVaR+7UA7x07IfmMUjKfQJtYaLZSSkeKPrtn+gDWOnVtLoLgS7RzClR68Om2D
x94E2BEQ6u+g4OsKJwJToHJ1W4xNGisr5zreYCerZB1JgQVVoAfj00a/cHooXlVL
EOTi1WrL4JoFcG5wrnBfJGVOWjUUX3dhwMrwg0tTLiWi71MtKRuu6jcO4jiYYiZl
QFGkT+cssKKN6IXZnMHKGQWpgc/uADYNGDKWe7J8vnPUlIDgyC4HGUn5U82gDe/m
qnmkru1k4zXttrYhlFt8ROaLOGeE8bTaQuKYhrl6tWHgrTKjicLye7FLgleDpfTo
qK/0Y58asqjFfyZMYKc9SgGs5NS1ACWNgbCdAuRw78RVe5UtDH+4Ryrr4RoigI3G
VoVaaAvsODpT6BE2lGqp6f+LwQEjuU8h+Y0+Mzo0bAXfc0HITM7bKRegaeAMjL7c
EXdovEcJwAB5Ej3e5xvD/LowoCxW5ASFUpiamzH3oT5sdhMHAvlvLfreTDut9Nkp
vVzm+ecUizHuNOfCjHSFr5r7+EpSYnA38kZXtV3311dMDNecL/dY7ipSGUKjAzzx
QdG7CcnpcekXUiEhAiNX1tiqTvH7sBLCesmdd6ZtqAKrZK9ygtiDEQUrP7mDwU23
fqpK77UGRmroNmtPKXpN3QULlKILjCr2mnsbJ480XG4VlX0u7Q2LOu7EJfLcDDgq
eTkIKuXOB0kgYmdk2NcMpl+5+YvFj4n7hymO8PfccMpexrzrPeTrqmB7r3AVFRla
JIrNMAf8sPib02aUq8IvdAyznrDNpugr793kdhj6uO7y9r3S776H9T42PX0nor/P
2Eur5psYhNIqlvXOjiQO62owa6vFtXuLQ7CCw0QJ0HZlprZNNbxIoEfk9bbtQCIW
PlNWdoJW98a/stLxll8E4I4TctNSNW8YVi1D41Sx5+FZvwDX+vHhcfd2kSx3L2UM
ZhrQWK7dkGjx9rWdvo3bSg8brR642Xsf+aB49xZ2BC2A92vRxciDX8u6y1MAq0t8
C9KB0yUtwWdTy168yfU6c8AQ+wv7CA8PGkXkr4maqsU7qZBh7G/604jQJOQv6v11
IZCj+ogEBp/4Ds8n6/b2MdMJnYZpDMakhKW8U0cxOg/GrzI3kHUX+qWO6Ppk2C83
YlDCx704SRAWDwfGNB1hBE73EbV0HYsCpw1PrFV4GqRuxGmrEBGGfVIilpPpGE9S
y0BV+hflOO/99+W7Yp4grVAouKlAcE6fyZ9E8CVVJbJ853FsOgY5e9T7sBszBWiD
6/QWvwAsFlcU1QgR7UDjrSE79SF3Rt3ktTbUUHhL+iRHvtFhAs3XMUxtIXkvTao7
/6psZW6nkN0xATUp+AbBs+ouUboxdMmhwk+92emFk1aXDjyuB5OAQEvEC0chN9Ki
3ti1M5Ye9W4IOZTz84em5GW6Upb4yA38gboij1F0CrZPmVEpwzhr7hHKUgJzMyz2
00pe34IwKNHDFm1ScCyk3tSa6l6hTjFoqhE4VPV7D3p5XpRzpZd2EaBXry71CkAR
8flcZhVoygeCi5kloPl0SxwTK5CSFvrCxAIequ4qNY7xMaTAgFvpRKx2AEMwe80v
8xN/9VTiodGqv6mOXL776ZZlYcFY2gxpraeuec0+5vc2i9ZPVXCaciyb57yaxCRk
SKxau61vdfex/PKfE/bHI/0g9Tf25x3pXfksoLir9GFt1KKjp/UddyF35ZUy/Rem
BH2SkUKueM53dD2s9GYdTu9KAbB0Fb+FjznCdmiXwpG7Yo+9Y3/WkiHHgWrnqCuo
Duhjg2nLstwMvKNZRxRZDUi0MLuKpZMwbOP4zQcnZ/+2aGlv3nStJ5vsKRtH5QpS
6JDAgovdQiE8cEUSLkutE1HPRjZX5XhrrH/wa6PuOtFGrgTNVPnXWpSjtzG6gOdl
C5o0xiwlhtBImhFdfrR9VvpBiHVebNFUCl4L7oWhAl5Os62spb/lTx+M65jQ0fFh
TEKtt8EsuT7MZckIUs+p68nxsNUJCYDj/aZq6PhZ4ze5174ElzSu0D3GAaysy/n6
nPV9iK+VO7EX6f0wq63dFz4femOi6fIcxnnMD7GY8iCcHHu3tLjcisiy6npxYuAP
OvTe43/zxudF4Dt25MZzp3As2FfxAjGcB9ql3gj/59nIXuJPchqr0nmvikdI+HjW
8mRhcjaozDghuaA9NNRewCdXgTc9bhe0g/pqxybK4QImJ59B0G7yME7Mcf0Of3WU
7CdC2OJX3vkgKrLVyRWOwACtDkrLMoA10sGJS8VTR5TYOYV1T48M8YD8EF9i6V/8
crMUPCTJuUQhSG3m3vjpdSTpku2E3Tq/IhO2qYGQly2IKcMX+Vwi98omyvh4NN30
1LTnSKTIU2L6wHCakVXUz9TlthGvRlhqAiTxRjzVWELNYLPj0PMWMygLVzvt0hKJ
GN1P6KbLH2oFNxMIyn0ChyE3I+CORyitPctWqAkQAAR/lm0UIpPH8aMBCJmcyAdn
Uc7iwDrOkiklPdLwDET4mWr/PCkLw/1F9urYgpMEgjn5r2hXh217/w7T+Bqgjvnp
XfF5R1dQ7wMmDe3Nec/SPF3Jn2BZuyhSeGVfzM/tObejc7LwMCD7uehH2R69MiHV
fhq2AbmKMPzEU2zpWgnCpq16UDm85QrVhkDANeBsJ4S3ihH7ZBtlzg6vycGR7pYr
/x3SydzW36jcYIejNjyYnmKsLEuoAbiOmSr4ExzAfropfwHb+9BJ6jEnzQpgTZJC
kx+J92faxswoInkl6Ldu3Y5+MNb1ISId5TBh+5hd7vNA2ZdJFm68kfSRGWe+nAfB
jEZniUHYl0/i5xkqBCSLBP+fXCHSVVqB7Rs25YnmjP1t7KFym1ulr0F9rD/eEi/R
GkCY60nfOiLkT0lVSYFT8CR8s4CgTqaTPkNJ1kRoGHFrbPLOVq4/7EWh6P0cpHBS
6NRyZp9GIEmWNoUsKHlrH/+BJPAuioM8/vAk+rpR72lUUmcmxPTcHXBierMc8cQu
F0GVVXfCE9QzSXDeLdox0+1Zi2aYMkRgsZgy2JMpJ079eXpLaZXv27QNr/M2m0qg
v7BxtocZ6KlopCyvNYrVRQXZ+J/I1JfDP1DYnj5SpFSYynmazcBpmpNV86KS6PRD
HXrOP7/pCliGM4HpfNKqb1lqpMqBVVTAB+H0dj0LJssxV95pnE66oH8nqZJnaazp
aWu83u2WzvUMcOD4f5GOBI6B0jJ9nfI4r6QczREY8waZCZPOy6tSE9UUEm0FJ6Ls
hVTjuGfU4ZLYOoC7kQb3SLJnyebCigvkveQXLHWkuED/mdm/k7ePx+4jnG7Kr29W
Yz1IgX5JTw0T/15m+jcwu1ILlW8RAC+nLtuRAYlBL1HZ7E1HBwB/QM3Pw15ELa6d
yh+PTnUypKdC6NKYYK/gVL99EekqYbM2EVisab/WKYORtIw+OjQ+OMQXPq+Pf2zc
LMGBXFnAOvTcpjzOxgxFvdaJv43TTlMNXJsqhwhROXSozKym37YNpRHbqnm4T4xn
TBKekPNVx1n1q11F8PPqXcxgJ8S1fDGCffnBoO51jWoLuZF0YB5i72wJUFVQdxpE
YS+npxnZOVwMC1zGqutvuN1Yi3jJmRdPAgnfMygUAEFqIGlmscpVAYqwcLtJ7vYX
/IHb27kFvSpa0kJ0rfirc2KE/RjDSSK9wpfBkVj5m/mmmtQSFMCy5yj8pbuZzwZR
wYsB5LaFF3Mo3+yYORVMOU4klghaH2ftNWExF4CAmRGaKZYM6+a/5ekHpNnGokl3
QQAo+FQ3/sOtETLRVOBCneawxZDQX9o5DCQp1VmyTTMAMDeI2W0DVeMW51PLg+IG
9SUJr6c++1e5lBTbWtlBaeRpMxkay1Xh6gSPLRqCl2OLwjiXL0etm6rjK9AgtoGu
BJ2xM1YkHjgGpFPHY26m3iJ0u2D2L0TjMQw8iZwirY8TRh+JHAhsPkDm1yG8rFbO
wQSFu81FnGun1p8LcCaD88RVvO9Tw+1YNXbVn5fJ8NA/iSylfUsDaCzsfElof52f
TK9jcn37DR6wSmLQRvo9QLZF04OH0GZWJhaXeM796MW4YQKD0CK5Oxotp9+1Fj19
ff80g0vvcxt799oSR7I02le8bdLsAmiRRalP2hSDbB3cGJjIZ1iRgSaxTQYKgkcj
Tja4FmYQb1L60W1CmkQRcpcVFrDbBLmM5Q3+ezMFq0Qq4l8acHTWvXMOCoAYDHFu
eTz24IYCRPpwlswEDOgy+ZF7ckP6FbdhU+xDAmMMTttErnYXZng+5fIAhnVushML
oYKEhg96+b7FBWHzGryTNOhuLXx7WYxGWe449rN/mxtH2X49r9yYO9fG/ykxjGcw
Q90tguQIgTheOL/4XPtP2j3wFJ04DE/riaJ6xKqNUaB0OwHT9rAW1I8y9NcfwS1T
0WS5G5zhmJP8LJCCoAah2rlPw475xmTCui3E/EruicaAIadnVSwIBmqWw+E1PIfX
fXaik6hT7CkNfDu51V69w/4hFhjKuQ0LKVbTZe2AAt150GIrcywpd4YRB83dunh6
Izettysrlro2/nJsOZiH5CQMn0uSQmCFDBqp0gQJ38y0FUGHMrlEuTVAUgmdfBHR
SSSTzcp1OvYUKqxLnRaf1he6l4Id8avTCaTfynoLIJz2+ZVZmjlJNf+YBmwiUTVZ
9+s7JHfaCmFiUbbYxJC2rP9NL181cbB1XGhkMOwfIbR2RU5z8ZJWMr5a6ycX5atO
8GzbGMdZFK8BYP6KMwvmDA==

`pragma protect end_protected
endmodule



module SB_RAM512x8NR (RDATA, RCLKN, RCLKE, RE, RADDR, WCLK, WCLKE, WE, WADDR, WDATA);
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Lattice Semiconductor Corporation"
`pragma protect author_info="Lattice Semiconductor Corporation"
`pragma protect encrypt_agent="Radiant encrypt_hdl"
`pragma protect encrypt_agent_info="Radiant encrypt_hdl Version 1.0"

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP15_1"
`pragma protect key_method="rsa"
`pragma protect key_block
bLj5GwB/YGBkTVvOc0ljUxu7i/SJvTvj8ulqWbVPwY+4jwyi2GWyJ741wSacSUdh
i8hFdRgNxrIqq6WDd4rDjnQ6ELO5J7xuy/y2ueJvnVXEuwgdndw3Cz8ErDogTNot
lYq1QLJHcMRydQxugwCdjtHbtGJXMZ8YShx4aIDgAxWeBt/KGIysP9gqUy5xKDL8
/hEO48+InN+mxJjm1ZhRJ5zMeWipdsM2StMs1o4fD4X9dSSNMmwdvHYnZMM8s+SR
k6nr4CLy4w9W6tbOk1pG696csl471mF6ZNTfC0cysnM1XgHSdWO+CeWGPRPpBNJv
8fc1N6dkDlFo8Jmc0Az4YQ==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
GNPdehrx+Jjt7jO6QLJ5UbvnT7kEIK3YaLT5WS96/9RxxIOxJWbbY9Q9fvS9kz6H
dgLUB4dJpI7bZgUnZmmYb3MtwlAi3ecNB+VJjoVE/3cZZyK5XQ6CnN9e9iPbCXrP
IgNEEfRVhf9t/Yx55TwXeqaQHimS9gsx8KDzT9j7mxGFuq47H5ORT21uXjJyqmJv
AXIjbJYTpBx4WgCq5pnH3swhrM1PievgLI6Y18BUAsHhZF0ddYsKAg+88uGYNah2
qG6aUjvb+r3xYpn/3d44SCZ7eLfNrNuhWdmSDUAoGo5xE8EjZhALEvfWsscI2zz5
Oyh5QVSayZAJVB9xKWAWSg==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-2"
`pragma protect key_method="rsa"
`pragma protect key_block
lVOv6VXTQr9MSG7I+NHVQ7AwRMHMhpGuq4OBoaRjytFYafq72dz+ugQET1GUCxmZ
Hk8n+pm9FIWClF3jIS1kEvLH8WOQDR99N+HRFXsqEBd2yRT5fqoan5cZLpmuwPkB
fY7/+INHeDY8DM6Db8Bblj0sFarcEM0O+NnczBIcBChM6k0LauDcZ2m5kEwOqVgo
RZC3vmNDd8DXg8COnWtyKa/xy/1KDfa/QzesWe5fqTqxee/8VMOgKe4VHmGvYFFV
CZkVAcEAvPAMtK66+iMbtGJE+61s2GMF8unNii086iRp3o0m2o0fITI8eKp4HbJ3
N1t+YrCBy5M1gTpVYuFyUw==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=128)
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect key_block
YOaeMxWkh1bAlcBdnU1zJgSKDuFNMBTPKJYJwgMAZyOPSQqBw28vo1AuV0Wg30X6
1RtewTyoZ9qZdytBs9in5HKWyx9eX+Lexnfs8cBQxXh64cWqdgBbGiRZlPtjaFZJ
gJig/ISanJzT9LCpxOolpmHsspT9+KS/epzYnQTbtvw=

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Aldec"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect key_method="rsa"
`pragma protect key_block
xyOR52S3+h1RPfKEX8OUg9Rvu7mIW6dNxmq/z5WH0ecxF8YfzcTYqL3LaOwquVg1
j88f/zXx0ZPG7oc+CI63Q+MXrSktctnaCqcLB8FaVRD8EOc0XscvRamJgB63wuOP
/8RkpwRJMydCwmaO1XW4hvsEabrQKHZLVWso8ejgC+v6yd8R0eTnpReDlBpaZsSf
tsgfCGvZbZ/K+nTCSFpbJ2fgg9kYuMzku3pByyinVDyK3L7na3D5GPLOwJpd2OZu
1Ygx5L3iQt++zgqNFTCo+qq2OiDS7rrIXdCD4zWL70ib9aJse1wZufP2U0uB+ECn
Iy8DRmxBl1Oknba3Nwqmjg==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect key_method="rsa"
`pragma protect key_block
AUzFT5aTagH3dZEFBs21JOICYhoBJyyk4kbSOex3NN3woEuNnIpt+a2wau6Gdu8T
9ao55E057JLxYF3OI2YzJrOtc19Y3sGmUfogTohvGpNLWBx7qFSzJdyk9Sq5JN26
qFgjoUys80tD0WyA0AXerVSKbMGC7h1jxDl25PnUTy5h2FeI/byI6QiCMER0ulhV
69mEkpDh/R1QKCI1KIZuI9L8GX1S/NfaJmJ47uDTDePIPGwbGmqR9mQMPFlY5SJa
PPh0xovI4l9rhlPtWBZAWHHiQf14Vcas96MEH/BDfBOdnKtrv7K2JraYtvUxmCZO
Dk+88D5xjAHcE6HCAANIlg==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Lattice Semiconductor"
`pragma protect key_keyname="LSCC_RADIANT_1"
`pragma protect key_method="rsa"
`pragma protect key_block
jvm64CxvgwdVASTQmIwlsLdc5eT2k1EZKMjKhyVH5x+B7jlL6lDtzJkBmInC0EVW
w4IMyH+Ls3WcUEEDWQAuYUWAGlJCAWHwigtWnsQLCBt6xVGRsgoji1yH34Or3gJI
SszTHjPEWRYN0S8OgPclmf5X8pR3uPzuKvtfWGJCI3mI6RZiikHGt9P8TtxJ6H+E
Hj5p5olEIkFrUwHhXnQA5Cd+Yp8Ph8w0CSE3VHTHtnnC79Ds/2GuOZyrfNsoLmG5
1QTGhI869WES3FPIW8k4ZVsWVO0zjETvruihbbThYfsut1DEivqGpD9uenLGGEbN
qgANq+7A4XhXfIxwQH6Kcg==

`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype="base64", line_length=64, bytes=4000)
`pragma protect data_block
IpxjQtkT10V8CGAntyVrmS306YFCUXBXNUwx5dDDihgHHa9N1BVUw1UZJvKbR2QC
bkuCf/skaUyj7EOboe2Pq7o6mbYVf/cJdYzRD8IEmeph1rKMCe2TbOfR3WtGerUp
QOMu4mr3akwoY+S8LL1/0fnJm0MMZg3wNrhQ8aqgv4vHYus3+5ejH6xJhYdAkN18
5UEOaEDq5VuC+xIXNZ+M/7cUs2nt6hUyWBbsvxLaJlll1AoerhHRRDDfM56GnZFh
SSIvWya3U28y7QJ6Sh+G/k90SRnd1Z4sM6aR0UnCYmIoEPhKBm7O/ictTdCcUH7Y
Q3ShA/sOFqUNfSJurzi9EdP95coUGPL2N277WtUgeg6UP2WyfiqObP4rFqy033ms
Hcz3acLOc3s1FiTPeEc6WDHRA1srTPG6KmYV3zAfRD4F+h6ioiT5icRqDSDk8Agv
QsM7xNPyuXbsGmz5W6lGWGay9ynCpU86j+lxjJEwQJjexMslJcgIHxz647u2mjGt
WHXZwiJne277g4Qv5UnoMGHUve9La/lJq9KmWX+WseB4bjJrGxNO8aEnr3i24Eu5
o2K/qZCGFTweo6PuCXHc+g5sk7wPfLjVQlvoHLAbtjIuNjivlKnE9hxtWXOTp1MD
VafnZtlWxk3GKsufpmMCvv4Vz7sITWPMsYae8UZGl4VhniYhem+nODHNeYjXQYSa
ETfPPylt4utlOG7Y/Pxu7Xf25l1zKCMRV6enFJJnpVZxJMoNGCLqHkGpiZ+JLm4J
90M7sgBDzPJjJOZDlos1wgf2Xt0cR0tqP9DVLPoPQYHaUZSp5skyobs9XzchtZye
Gy61KMVvtdUTahbmTcmLYn+ojH8qVBmEJ9GW0NwWca2O+bKsYuH83wh/Fhofk/+N
BX5BlOrctaAWDsA0hVIXg6DOqUtFlUlSn3NwfhSc/EUyGTKt08AV21QfVJ+Fv/Ti
pgAMnwtsptF9xsju6ImMJ1A3yOroMsxNUa7/xqLS+CMfODHDOCqo+xYS2UJP+664
GbdI50F4XgbT8AbzPTlCYs+wYQBwmNO/N+Lj/m+j97+dVKlp4rvHYTAv2wuCuEE+
XK9cuf58zs3YChzAjBOKJcrivQJPbuIOqF4guprvB92MKzlYxMjdTLC3a7mGXaSQ
pHqPIOJYXlLTAQA8UFqzb8O40xzuUQEacvIWTjnPLE/DhV1L4NUhcDX4JUGPSIbw
9aijn7SuuzufdPCr3MmDNI4E7DTNhaVNnbtPV/WXMl+GGQTnwvHjnVPamXSdxe+N
X4uEOJteg0wlMJ93dD/xT8mhRNAVTQxgL0KZ1+UpFbFcw5/MR4BzFYOmfzlITogZ
azqDFMF+d8VsBxkbMTHdraR52ABrcNenrd5XJP78GYXbQfwN5l5sXbZgrHlzPUw0
TBBavDKrbTkRdf9lbn5/xdA4qngpKevvT7iti1QDQgCIxfXCml9PTIKlGIEZTHqJ
udFxQ9OBMGX0fGfliFE0qf6bhbY+AsGxEaicPtA/gj8+jXuicddvUeIolnUzltJx
fgp471+cTfv3cf9Qz3hF2xOLIBHU3i1Y+lvwlsVHcOETLArOCBm63nH53Kdpwtu3
Kvej45JTstSXtNt/oIgTvTmyvlpxAYyb6DVKwgztcAHb6UUS7gkEiDwAnW98iRO7
ocKxklnJ0x+HLzyOY5RcCs2G8y2gMEOy7g8PAVPKS1FLrkZwhnkntVdgTpsC+oWh
gYeBb9WBrNQ1PAZ3WNV1T0M307HAOnrUuYgMx9IJkQ+k5euWH6Fhh5nUB7BvJ1hE
N85qZrUiO8yFGo5tWQQ04PlDlRrZg3eqz7tUEqExpRjNDEF3LpK/8N2CrOb9cCp6
dhcYwKBmsp1gUM4ES+mS0yjhP1lFt8y7LvRWPDbEodz6CElHSXNp4oN1CAK5mHcV
46tskJf8ptlQ7NYpnq/REJtpPXinXQxQXq0tSSwXDhFH5Bu6ngy8Bw90cCw0+Hvo
wbTSy4zLUpauyHIRT/5X/fS5tgPGfJE6fX6v+YDPOkfyV0c1OiFHb0IjmSNY6/6v
9J/DqGWFH+hMvzdRfesRoKRt8hqT61XXqjN5tRMs2x3YM4pZBzeJndzDfazc3wmg
6TXSU+M1rEsx6qnB9SEVeVyyjWMvn7qEXzkoPonWTHVvdzSiQU/YarJaVZdeP14R
pIiV5u7ZqpQwDvtLjlgqDdRq4j162iYP1YfEnBuZE5eF2K0qNmNHv0iKKXFNdHP+
RNknY/kCFsp3uIFX2k8Wg0/5SntcbJfLYNMBCdeKZNkCVLL/kf9KeEEG/tWRUDGr
lcfGzC36L85UWK6KPxIuWsrPXPZOTTBGlKAI5VHzW1qUSGgqUGjbPx02jMNEyk33
/Ii4XpE9MbCzY+N3Qk7sfPYnv0qnWbNWxSyPII6GH+HHdkBuMsr8qoUGYASoWpfW
lEQ/AMDOM6UiJGaX3tj6ONQWqnkf1DF6e/b3ujYe9GbwXw0Kd84nTrY77AV1hUaL
L/asXUTcdSWvubJYR5/yjs91wOXYpidf4AQoHMFBTT+KAqoygyZBBxPRYmVqFNkK
OADrrXPaooK2G0kIg7mbYpZifEmzQl3ffvUc7WIign546Xstn3w9Mio9hQBAua/g
cK/d6kbjOj21vgaB7qy+thxoU7LD+F7Qe0nwU2QusHUVSw66osWFXJjkSKjwVINR
4GfVNNTWbbjWpUwf8acC5v72yY3yM94IqDzBuoPzCAwvcoaN3z8qqyRrO6b+ou8u
DKG12UtAY1X4T7/+cpybfxnVViX4ujhOgkv3zJuQhIX4LVtPVesOoLJD2GRIghyb
c1+svZewORNuiOOj0a9thEuifZ5+omG3DLuhCEyRJkmTbtEk0CwCUSgqWWK+/MNq
yozBFIAD4WfV+liIyYElyjL+uqWBF0twKIeF/3c5lejl6fyqKCJwi6AIHwknT7m/
jkJPHjkAGafR5Y6RQvXm/Cow0VAKredADw4DcGKhcKiK6xucbNnSQcc+G4CQuzQm
w+KSdmWwuIvM1C9qZddtJODWJt08wEJhznjz2R9MAQg5pl4f2QIXIActkxgPmPgD
hk9KcxZO1CLTq/3d4Pg1M/4oJ8buCFzUkoTS8RT0b7RWXpzS0p9q9COZg9u2dosy
L8Y+JrYm9bX0t7IxlEOWtgRSnjjJSeWt/OanwWA0QghLbh+AzvyhpkuZEZrXwPtn
U4OzpNhK4Ti7X3mkVts85CMMfxr0avMlYfh5sDs7kYooDFDFmUWLq7WTXe81a/oW
A3hj/MkV0HnsgNSYOaTDtqbjBzU9RsLawTQNV/BYJEwZC6ANe0+K9d+wQXjJn+Ud
ru3aAmWKXwinFgUqumGC4fVTApVu12knd5Taat39Gy2Q0fwLO3/h/w03OMk2b3Z/
9Tq5V+N9U1ilIx0Mu6nY9FgPt5qSJoMFIZJxDnxvGp6wAaA954EcGkjm3UpprOJ+
azTbeLYT/+ftEQVCvRd7sNzAo987eRgTTuQSap7ZPAycPTa3IYg2e6DpBeKt4egE
bwCYamj2+dsFTRRHoN+037I3vH+mc7tZI3YMDUYicEyfr1TjCQ2i/xcpLbisg9UL
KkjBnhfJPp31eUzUvpbBpC6xXk2xIDFBYk0ls4gWJHfRgp0qd8y/28I1SAY6Kl3C
KW4F7FR57a5Z8+8ZZVtzOUTWA2c8DeKJdQB9RnZ2FGb+CCWkWtl2VFIRScCyt31N
BFCTZinDdk3MOzL++7wrmQV+2q8WmIgBJC2SjjKxMbCl69ni+IJkS7iru3ZutyRk
GnA3eXkn8bznjTp2ZhWPBi6fOQXnJcR/l2qeBpBquEXF36coZEkP3pM9MUz/wExf
VRmc9ckOJDe5mv3HLaJnpDv26r3DocwacHus8dgOglZP5AM8x12ciFLdK7CM0ffY
FV2ii1XcJggTmytoGOQyVLmbXSiUyx/BFhtcfB7xFWg+no2wqkQUE0QmBsCSEGj+
rY48Lt6wucvaBtj5i0vzLYU3oYSOBrezi7ueQBjjXf7idqGXayGbkwYm2h+k4FSt
T+cWvd7W3hfbSDaOJikdY8I/6E4QWE88iY+HT/Mts22GYFXU/2DHKeXSTuj+Od6Q
EB9hHGmkdV4uobcL9aHaYUnNJv9n3yPCLJVGcOdUwxkxrXVSlFxT2EgBx1031VBn
n/NwXMOAL9fXzulfSx7PLJJ8O7UXGSSznC2JJ8KcHE6Qf5GgoV0IcRTg3pPw9gZw
F9JGiv/ZCgTAGTAFI0lH8ae+h01dBQxihZM1u8H/YSj/Bjtw2Gowq7mCBCnPeJMT
xFjIOPeHbaQplrVeMzVJ+OxVDhR8Ph7p8U+JRZGhKCDT0kieYadf5rZWXgBNcpo7
W7QMM7a7SOjrd3UFHQun15B0Cz9Pn1px+0olSqffL8tIzsjMqqFZcWZTJSpGQLAL
r91JRJyd6aQibU53mWrzM7+j/TD3J3WQnnFfOULA0tayu8vA4H24pC6LcmVSPLTE
xFx4YKXpozsQJ4WcHBMhBMe/IG2Z+pT1mPhYsWvsSNCQ/v+knc2jwVz8Ju1pQC/7
swDl2KMEWZKXZ3JORTMuJVeMwO3g7A6SHHjOP7sr4jctl+F1u00+qx++aam9hK+j
84wk17CNZ7WGVEOtzDdsuj5NVe0KftNTDsLvObWXO/06UJIvQDHPo+8KDRtc0Oui
emVZuytqQp4HUBLpJ0+1RvqOURGyzrT/w/HYub78mK7FRuwJxSvtWGGK/Ni/ZSwh
Gckf8HbXqni932kmiJJ8+ZETOOvJ0CaDZgtKjttzTtrGZrZ36190w6OQ+R2HvdZl
HeU66ciXKCQKLTVg0JVUEmd6blCMRoi2WX1GIuT5wnFX7O00+Eo32EJwR61h2k7K
ZCsDVmV14P/fVkRTZ/dkcWUxLbc1fkIVsMu/RBPIoDEjemZ84Bw5XBkuWvz4zspg
DUoCAWh3o4kC4lKARLDNNMFJ40KgUd09UeOGOM9CBDYniqsAeNio0TFqmG0WBPYb
IKMQvU45UYMuC7WIUVzx0/iRP31lVcBEU/dvR9H5eKghN9s447cfhabI96Z3gxrj
8oGLRtJXMBEPlshAkNYCyHW/djVg6wnN91lSJ5daMC/GuHYJ/vcOEmZP2MzhLKGr
OgmGhliaVDJOEtyixfId1ZncjvWI15ly42qrIS0OVrdoxHPRFCrT3fwcnJh4T2Sn
EqkrsNyGSNInkDMTI7OxkwUfv+ZSBd5RvI/EklZyZGIhS/W3KcO4eyHiTzQ/JyO7
Ii5Rn51vcXWCrrKtsz9xaK6ORv/FkAKE1tA8TNJwnaaJrqLDSFcabWoQmDCuY4+b
ygj+ZcEOzbT3ARks0kCuIQ==

`pragma protect end_protected
endmodule



module SB_RAM512x8NW (RDATA, RCLK, RCLKE, RE, RADDR, WCLKN, WCLKE, WE, WADDR, WDATA);
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Lattice Semiconductor Corporation"
`pragma protect author_info="Lattice Semiconductor Corporation"
`pragma protect encrypt_agent="Radiant encrypt_hdl"
`pragma protect encrypt_agent_info="Radiant encrypt_hdl Version 1.0"

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP15_1"
`pragma protect key_method="rsa"
`pragma protect key_block
ecgiXXmhflspGVWk3zTGrNznm1/aJMLEsGuiD9PctoHXQ0jbsyYujtvnwXKWYJVu
sEHjlCrsqX6z1N4yMVvuVywieRDhEtJFQAAorpU0jsSNU8Q/9nukvasRfXtV9YMw
Hs0+0SrXQdSu5esNixhwga8qJQMqkQBrfRdv8+zYeesO+QzXNgWHbW5lcNflgBTo
ziOlUawyU9XHRNO/W7ExeYMaSnSWEI46WAS0x9iCUCWNJK02D8von8zkLqdQzwBh
GoJWY7uvtLuCVrN4WbloOYe5ybsWcItWaMV7J+GWaM9YSbkLgegSNept2GgjN97q
WgfEn9yL9OfpI5a3oMiS9w==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
xlQKnhwSmtqKOnfKFU+z8/i3weyxx/OI1SBibWpN9882LifrSzLaWNZ4b/7h0L5W
Y4juN+65kTVHWM5r0Uq6omcPoKUonAS+UEvjLuEGALm/XPBLHxWzcRtupf4ojDaA
uJ4gdNP6EMb0nZv3NBqrSktkIUVA9FhSUgiNnA+1JMV/awjiGsHyXcHm89sxLvfl
pxhYNaqqbC8vD2FWi4YE7qf2Osts9rvVtXOlOlFtNfWWt4VqgaukVvk2B8i6BjL+
9WY2KbCb22d46OltN7JFzMLJ00wqHcNAUk1fG7RDlfaLkTLV1A9Kw569cIIMQDAQ
v4n5zZN1UvbcVwwAW8D5vA==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-2"
`pragma protect key_method="rsa"
`pragma protect key_block
eGdBlWpALdeuIabjDhIOUar8pWpUPqC6LKa64lLE1SFjQHeDsmHAVrQ2C9DtFEG/
QRmhmbxplC0BQ3PlMysNoONpPKLxc7GFfsFoRJ2UG9HXuTXz6bwOFHD9oQVNBth0
iWO8zCU8b8eBqywWgOkUtFiZVmMmK/k+K2UNxrFCXaq0KP7uisX6dDdhnQDWZpRi
bpZcHVbSF03oRBh93zDWBBCUJ8QfwEJQtbWX2fFCeWpK6LDdfrFNfuby1Fh/ZzSJ
Avf3nttHgyCHYcxLuJGPwk2HB4YXIiknzgzR6vdN9JSRuwedMlhGPag2KiY/mM+Z
txarQneUgcu9DELyh6NeGA==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=128)
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect key_block
Au0kFWiBOgDkk1n0NTRtUaRfHpZH5J1elYQO9dsBoHsEAJp2QaRzX23K0JWeNJ7m
QlSrdpqrktudzMXF1PchaIys/lQ6iUWn5y5P0HRaAW4jFW5efkVcb1nR/PkaUYYX
O44gcME8To45Z2gd7nvkfQ8wxWFtxI5x9jZF0gBiJng=

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Aldec"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect key_method="rsa"
`pragma protect key_block
Eyy0WECICUHShV6PBw+0R3x+0vkCjLwHFB0J15acPqKrta6lwHpWbZLGn1nCrk5B
2JNLRQFhM2stBxAZYAHCkAu7RpI1WLp3+TX23iaMm5JuglB4+hpIicZ6ITWD3GH0
ws9bq/ut1c5AUKjqwKekp6PS8bzQyXoIKl+dilKZG9s/4buLdKVuv1WMBiSBQQq8
0S6KakDJ4P2UFtt+RDrjs0NUfY7rEeLCluOCrTKEXzsx8BOXWCmboG6PAvGCxJR/
mpDsLS4Nv8XPMuchJEO6p4FQkLAYZNQE++sN4aUZYOad2DmHgi0HiqC1iAYsqvT9
Rxvc2yb4UCrbZMQZM0C2UA==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect key_method="rsa"
`pragma protect key_block
B03lv9HoAajUMimtW9qOTZ77B/MflEULTqjIeo8mVNjB12MN/hkGWyUNiunmM3Yy
nPmQ0mjXS7tyD9y9+U/KL16M7AkfIx8eN4d+el3Xv0HqJ34jwP6gLUATDOYbyO1x
Ubz8QAxTa68yjSbaoeZgMelSjyuF325nn184CYt+pmYGKIkLAkCYgMCRyHkEZJSu
rbcNqepBAwoliV5A9jjbdxPYLoVKDOeQr5sAmo8K6KzV1ehHEEtbeqnraLg5fF4N
D0xus9wSu49JlzVEetUKa+qGfcAU+DScXD4kdXScopOu1tGg6wLoxVs2xbZGF+1e
MOXg695UlRiWCZITYsklOw==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Lattice Semiconductor"
`pragma protect key_keyname="LSCC_RADIANT_1"
`pragma protect key_method="rsa"
`pragma protect key_block
J9WEGcikoFVrXbqB781a63BtWy7heeiTe0OdSv4TfNda9nNqTNih97WXa1qrfSnn
A/tcPqlyt1edwP6wslEVOWEJmMdPKeDAKS2Cu2s8ctHDHnVUgRETvMaf5sHLp/kS
dsrBtQBIz3WVnZy5czZRdPLeH6rMrdmrO9MOq4GKJNb8JrRd7TEJgmxJdX6B0Ikb
Nf1Vxf0kgrqsDknpwnnJHi8MnJU7uf7pwyA//NCyyiJ/6cxiVPnz+Q7ueWjim2a9
Av7g2IbkRyXBKJLWJkW6huVUPJtHMBYcOIZIskvsdVDB8SCG9lm1qED8Wj8OTbyV
em3Jtm6PzL5bldwKyG7sIQ==

`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype="base64", line_length=64, bytes=4000)
`pragma protect data_block
lDaT5A9FIYJYLajbjP4lkoW/ldBGlSCrmhVDUOhtfaJXEAwfzBr4y/f4uXZz4Bh5
3aCiIaHJprIZOK4MV0kteyKeRNDNn/9CKwvO9MpqqSC9MaerKX0Y0QZeXK9+M7J8
ciG5k8udulidLNfSTiWQpUhTfpuo+G7sNnwTfMtinFlE1/8kUa5gcDnsDNTV8F89
HM/yx4gLv8uOpSTrcBsE2Go0lCtMtxV1u3l2kN/xs3AUMeJoRyC90IC7m7XVU1Nn
WsB1fzvZRfXv74Q0z2alwIS0UBnJxh9ZuRlTRH/undj5/EphfGq0o74aQIxxKFVr
SRFp80OJGL0n8fW9ehFzzeprCf4ClaAvg57bsAxJYOl1axLr8l5NtpfmYu4DWTfn
i6Qa+I+oQAHGxw5MySwWwr6rwuudYcPguzXnIX9vln+NXO83KCALY6AzReJdTOAK
fPDq2Ktl822nU6r/1bW7Qb9/6yUp+0fAVajZ4jZEW6trI670qvOlUDYXtOwRYz0Q
i7dCeIzJZj1qULFkFwgbMO8+T77R0HI1b9uyM8tf9sziwUdB6p6/RhHjGSdhnKcR
kLCw/o+ODGeGySaYQh4PEZToOZpSHSVO/m47qn4V5J4IETOX99MBpvgVs9v/uxbZ
Mw3B7bpZ+OzlAcGzuZdJddzcAN3HWCLnGQ+YFjUWp9xNjG3T2ZM0J4WoR9jYRZMW
+z8FGd/g+VVOi1hDryl5wXgX7oD4u5YBazYO3R5bPsJuwDB9+CGuoY3ZnhAT2lxG
Hy+9ig9udOgm7lpbr2Z2PuJS89qRqNW2E/0TUu6Vjtpgn35regMXa03JqtPOeTV0
+cRl9umNcg/5PWMLuPHTSCbogcUY/51EPAd151bKqIfAIqdQYysOc6D3/HB104JT
I3CduGvRO6dvkDjSOXhfFXBeDh40B1P1w0Yb+qePVJlLJyCnSm9RBvkPDtnaQjU0
eTTzaLqOAgzn+mjf74f7Jvgyb576L/rrXj838M69RzkJvWZISJNu7LYj7m8MfNtD
qEC+WSiJG4kyVq6Q47rLf96BYB9fSJMXKBzwOjH9EkNj6I9tNkzTrs1jjh4f1BR0
GQF6y1IecC3Ap1K3put5OQj2Gs3m5DARyslE3m4xCOGTTBeHxcAroRvJaN7AG3LL
g7OslKWrN4yu5UPMzGDp/Y1EYfEZiK7+bzBSU9ERbJFLR3zEnDeqhob1lpjvQ/6G
lBFj8jLSvE7pklrkm337mJdUpOIxOwcmLAVagQbmR2dicwa02EsaPa9JSTqsSJ0M
ZJWHg0atQHMuiyiyzo8d6AqkIX8WzAbFg5rkKGh4fJw6bjKej+ksTFGZPt925ivd
TmvSlNGhtiJH8EU9q6BrDOyIJijEXXfXm+1b550+JF9vAFzUbLcoFxbyVFip+sz9
AaCyaSxxMpwPSTddLZ4QV8Vm5YjSDMFFEtWsuEqRpywSMi/MAdTgi4cLEdcvMeYg
iRDIUuXPe8UTBZCG9MN+jOZ6YaCV4mLlDz9QUhI7QqeZP56tQjS2DIMYnRMBgteW
vKtegjfQtKRwQxPFiCWTkPCBjBfxdcNvPYziQGQxJGgIJtFZ2SowUV8B6nVrtGwM
4bCo3OQ6i7j8i9gp8pTrJjZv2Pl+Uc60rKX2IV4x5l+crUkhZV6tG/jrZqlVc8nL
fpCJldiTegt8J7nf7pZWpgBt2FFM6KxAnxxPrpa3m6gnc9NJG37A0S3Jls734Xe/
EEHGTWkCBQeD5soCIPaFThWOSw/LSjgHRlr1vDH42EnqDmH/c80ArSGktMuH0i6Q
OEpaUpVSQD/ZaSiaiswPhXIkjJ9/CEa/pC8OP84OMEdwLJOXmXbFoFc8uxn+mQ6P
UIknB2xtrJr6FckLfc5q2ZSNHa6wdEEPKrotBXfwoJXdJGELKEFIH5kynWivMzZx
WzZqOSfFa6GDDHKtEQo8e5hUxnxgJ6P6vjKPqiMGf5YKVsfFkThQ+zF8D7TcC27J
/palkYo8rIpeWUfP9NYFGghr1EHrKyMCCwGGUkukf+Z7dCWDwCWt8SKhXJo1yrot
FvjJ7Wf2mICGR+EYRgf6xMtftL0mEQb03CBVTTlrJIzaGw8ZxnJGvjk2Y7QzU2yq
N3JP7dP1RPYnKOnXx2qZcGeAkvXCyEBAl/41arRQTl9eVys8Ey4uM+R9Fmv4xyrU
hlWQbs8QrwdZK1KYoayvafSZUvwah9e26YY9NteLTDnLYrp6lt6F+hn1AGirtrnO
/CPDLuXJuzjGBV4YNnPMzST9qrBzO/PVguk7/0pxR0BFxnG34FcX24HwM6+xHVAm
Bc3XXWmxBfY5db/zIozqBi/Xy3HaM94HtzvgKHjFcJhIZl4b4I9a+5b0aHnOVXW0
Lxzb/FDPfUhJsQQwE3AwP9fETVg82WGNvJHbZsX9H4Hauborfwi8K6lpzRsDq7T/
nS5UGRnTUPdP0DbuaNMUlyT10Fzhg3f7R7gAMIeNl2aVghYC86w7FF0zP99i4aPF
/sxCeYd9Jrb39uSqAGdBihjhPoqhBBn8/5HzSvKv1WTrE54J2sQs7j5Qfi1AJfVS
IcoIZg/T8belk/UlYq6HMv+PF87gBpeAWSIs8xUwcbHuVJIvKGrLBZ0X1Fe/EAl4
ZA7JnGeS32O83WOfYqWDdedMKegC5q03/jpgipZkSfcdLcf+OLb7K9eZjkMuDrEw
740i7/iFfUttW66ESv17/Rcj3K244/Br8kGwBAUuAXdQblkLT617oJTj1CySkDFn
1ClTnERuogli4Kou6kS0ztP2smjFkiY0fRAI49BZnxJjgjKSpoo29fT0dEsDFY+u
UJHr27kQjleVj8l2Lhg0nWfRGX8gmFrPASbAmxmJSiwrNaZpYACrfESsegWocWRp
4PWQ3AlcyYWqUlDIBai8tSEXfZ80FXusTRrQa84dxHdl+l/Gpr/UftaBBsAZQckh
stNfKcJ4VBKOSIUlhMW+Yauxj6fwWtbqLxqYB++XMS6g8tN4fRPX1Ld7g4yg5xj9
pdKs9kQKz02+yN4gDgJwzsXwE5ZjrNeXzTEjfMBibwxDDBTozJV1nNz6W+C5qfVH
w9iMMtZk8vtQF0/BQ3pBnDtdLn3djnpW9qr0G3y4QQoX3VdBGzkUvgRbj6w6hm0U
9O3Lrwr+Atm5fG3tXNQeMNV0OllL/+PHssJs08E9qq4KkBuUb76O1AjOY4JBrsug
8vsF2HTyyTOosAwa961PYk6wm3LC9U2qJTCBhtoLjjnZCk6T1C4+fwxNNVhKN+pY
a3xZQBhP1B0PIh9FRgeDh2+TeQQ8pA2EOJJ4OqQpHj9TzSi3SGka2nIFA5/eI/qe
lHAf/CdyRCQE4UwT4chtrtXsQrfDLAscdUUU31LXybP/w0HqSSER+jfFJkIY5AUc
ijOPNzg/bvZxIFfj39G9ERm+EpK5Sgd2hKBftNoJCWwBurwuNL9RW9wuxjW/5isP
DXLZs2Cov0hN/4a0t0N5wNG/e7/cy6MX8bvcLqMttvSG7AE3iroRMafCFAMVtipD
dPZYEDNpBc3dsdmvjWbL6INUBRyEhYmX83758TAQK+Vf6lGBYSthIoFPFvq9CRRa
1OW1VRCYBB1Z06yk+suYMoWMFHZPgSgyGCWwiUlv37CRsr7cvLEMUoCXe1fPZPQ0
o3/THNpCy5S040rFrnxT1VK+CvZV76Sq9w/xmgG4L9ahp/uRN/lmDm+2sJBM+lm9
C4DxB3eKzka8SWkxeqWIJeyc7HAvElZlpwncMqnWvegF3VzC6FbyzJrghYHnGc7R
imEe6Qqu5jNmfgkwgwfZQe3SDPB6GjO/aRjieL1xzVpgt0Gg0Ijx5VdWhmZt6rqx
rox3QAK5RM48t2oD/qrO4vmnHfr+wzddpH6dJxVbk466+HwZUbRFvy+SQRLsttCW
qn+lPOo0h8CO6WhZG6bSJo3L2aKLyOlOdlE/rQ/BMYhYzXzmhcJnOMtX4HP4Hvf7
92zef9OGqMHgymYVT1A4wyG3csJXEpzWSO1IdTC7PE1s4dRzHM2BAto0kc6oaOj+
hBBTYdjHsWqJAR5WOrColYa9UQ3BUdHiVeeIiGz14G6p9912ikbWzy8GcIpU2PuJ
yI8/y6gteKziKlKrs7rPEa0in3/EjNlkMN44eLUhFtvWA7tNPzu2sADZzY8kgNd6
DbNwKafdShBb8GzlX1vKq607ye61paPlhy5bFfkz+MU8Au1s7S9yp4AZE1o5TXn4
dKu2mVJuL61zOsMlb+Pt+3osqo9jWBPytzu9F2L9dzVd9Ie2278d3Qg0ldlEh6cs
md++gbFbqb5rCc0N/fxL+PbtmG4b/bS+Z/vx/eYAlqwAWQa5+cLa3pCe7ihyoKuX
gABhOTUbBieOMOhFlBBx9RzMmlwCvxs0NP/erEX4Jrgif9knQYo/gtfyFWLhNWBI
4xRu2G0PAY/8XGpafIpx7g8Uo9SY9yYUzAkeRMOy7rPj7PY2bL082MV72hnr7A+P
mFx9LpTfXDpOwc2oExa7PMhYcdAk6lfV1CXNAFMm5Ys7gm9e8aRD/kA0koJTqjlv
pwy5hgcfgVDXZy0I5r6XJ93nQ9BBNA5J7mR7KEBZrGTp1R+h3IFfW0xRCwqjf5Rc
k0YHf361Z5+f6cwXD/f532ZgLT7cymPF1fUUDIdihVOwJShg3fWHoFdxcBbOtKEp
CukFqW1ZUejigBo5qYORecbOtw6+CEubCRu7MfOIKulIw4lu3MExLlm8xVprN1Tu
25Rp7zE2acs01Fc3lZcBXGWw55zqaKbM5APuDx4KyWeIAv2TarJFj7tQ+3n6hRA0
8XsDyhSEnj3HsB5bZsrymiPQQZrsT6NXU4cpslucD/8jcbGaeacXcbldj5uEy3Kh
FmX+y7HlJnD2yCYD77+ONrDpQw1e5SsRttge3C+HCYlaHPdxeGmpUCkqSh7Fygox
K4snFMQnUzFccZoQklc/IiZ+tKDCpPPP1kGDNQA4EAqJcGr2zDs/0y0wtVLr+5M/
HiKSK2yJ/sypK38KJ8T8nCFSRMfDQIYmbyxpEyB3qriMzRmVlnHctctRddyRCV7F
3faFE9eN44SQ1F1tu3jOxfkFzja+g8QqkVyfAoqubbLTuGndlaczLDWI1RYh9HS2
F6BG96tt3QQTPmNMtUFam1FpgKC6rtEm1h85gM6j/bSFuGyUixhRFd9mVUZScAnX
RbGd7ejgdygAbPCWEfH3vbr3NJYc2oqnFw3AaT6Sl29K1848L0snP4+Z9uJBa0Tj
ur3/XJ8vbhETaahEhsDtRbSUVBzF5sSB1ksqgtSGQD2RBRo3C2C4Oeh/pp+g7B0z
3w0coBj0KE4Lx4F6SMF0rw==

`pragma protect end_protected
endmodule



module SB_RAM512x8 (RDATA, RCLK, RCLKE, RE, RADDR, WCLK, WCLKE, WE, WADDR, WDATA);
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Lattice Semiconductor Corporation"
`pragma protect author_info="Lattice Semiconductor Corporation"
`pragma protect encrypt_agent="Radiant encrypt_hdl"
`pragma protect encrypt_agent_info="Radiant encrypt_hdl Version 1.0"

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP15_1"
`pragma protect key_method="rsa"
`pragma protect key_block
O+gB3EBSgY7QbcgvUyQThPJLCWgnCatAspajx+IEnKM9oIaqiCo0zVF8LP0WiQGV
VOP1NHWMA50L8BK02RVFeCx4dNW3kG6yX0qVcrDC8Chi7idDm7at4qJQPU+VPpck
J1lRkxWZws+t9q9kn1eswtWemzKQm1nAqHVoN/eRlEOyc+pJpPesI5f1bhle2UTX
Ph8rV8QmOJR1+AMEnbOWEjamrllyyznd6bGzXxZzeW1cB96oLIVds+hciv++WROz
89Rohlc9jlQyx3Bvg3/YMgzCsRALlNNsRwRlvzmGMZW1aW8JG01ORYpgUCWRjfP4
7yL2v/H81KQwUbIFQAnT7w==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Synplicity"
`pragma protect key_keyname="SYNP05_001"
`pragma protect key_method="rsa"
`pragma protect key_block
bPe/qscTKi9lh8XbZYzuFwCfKEwr81sa4PS/KUaLm3iFXonbit11SUawncxSfFn/
kxv9Fbk+5uFGNmEq8vbJdvlctktlJSmF/9FOGZp2WJcSpbMrem6v6PeNWDgDWFso
XZrRyv5mtaJjJKyVrxa7Hw+XBgss1WMQHn31a2eeh7L48wZeN/zPcJ3hOkx733zv
yyqnYc+bo6gh5hzcc6z1Jsl0FXgmxmyxKWLFVuaPuz5/addfHUhi1Hfr8vGfosbR
7SrR78R6m9MjROIFA+BdJ3vlPWxzQH1bBvPeOj8j5+JTL+oRqok4h9ocEyRg2L7e
oRbWkwSInMPcQ6KQFOmyuA==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-2"
`pragma protect key_method="rsa"
`pragma protect key_block
ESpY/xrLCOcxprktpstRVJW07Pe5SU3nAWyUOFZ+2pD1ayREX+v2jib4TslFp8t2
JCarefxsORCFaiHc7Tx3LXc5zulaFfWnvsDE/S943D6DNq+WM1nVFm1fxXBFIbv/
ZYwg931a1JnTFTrHUHogFy594Hik7SmOBhnMsCtfQF41Lzu78DJPzfncg3SQjcCR
aA5FdSx9u0PWuoAqN1VQE8fGNGJkkJD486HSpgmtnEoCTYI+f0DE0rSpX6uuZqDr
pwu6+cTzqJ2bWnXB284BQHJk0yGRYzqV03+IdTK56RmsotH/XPUMnzPYcURoVQEn
Phh56Kd26Xa2xUQPRHfxTg==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=128)
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect key_block
CYj44BTErcRl6NtpxZb088CAiNPfPj8Ll2fBIG8rlePhp1DSXjn9FXopfNmoSLI9
xawJCs7YI7NDLieord/TcZNpKL5Ol11EprFguKqINI5uaaN8567OemabK0yl880r
vngNRVuzIHnWBQAuWqqK3CDpuI0QQJLu/XTkPRCrbso=

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Aldec"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect key_method="rsa"
`pragma protect key_block
sUpaBcC/5Vo765fTCntYtvVY8Gw+HpHvl5eILFTd4jp5xvbod43z6cf5KP7Y+iVe
GHk8mnO589T3MuxdYNwflrYxCtDzpQN770DLk8uMqOqfZyhsaIj/zAIV7qurtRUz
lINDfLZ17+TDwdNOmvXIglu381pFYbxpf7fA+qlusEfO9//kATyqBBkxBAB/DGLI
yt16o9r/CiLoprL+1QpWxcL5u0Q6xXVG3GFp10UQBwnMRwW7RplfWSAniQO9t9tM
UeWj8kVKypkQ3gdseR/VSSc4K3MdRj1VjzlsavTt66PNhGy/dwX61gy/uEcVdpd5
apdTx9t4iC7lUGve38yaAA==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect key_method="rsa"
`pragma protect key_block
RX0+ol0Mv4VxvZFONisbr7ogibnyHBlTi4qjkVL5gF/lreShPEpWuupHY20eWUGg
Oqg243Zocujwj/1lBnQ/JX/HqVx9uo3gfEY1fy1XA1wEamFlPNkZVdhoAuFB+h6/
4YGDIH3ogrVxq5wolc8DzvI6jvjkRnU6bzQPWBLCSwi8sam9c9UuoHxFYZUMOK90
yGA+tdwcjCxbnnLtIJs5xAVoDwoi2bK6QsBze0dQdunD6LOhUeJj59s9GiWZY3bP
IN7/Dia/06tHhEOI0KPWZgoh2imf7CIzWJAWSKrqgnkY07ZVaNXZQ0++5C6VP44k
hYOP0pSEANEBGBiwpIRTuA==

`pragma protect encoding=(enctype="base64", line_length=64, bytes=256)
`pragma protect key_keyowner="Lattice Semiconductor"
`pragma protect key_keyname="LSCC_RADIANT_1"
`pragma protect key_method="rsa"
`pragma protect key_block
ygcPOIHAsH5GHUEaXBNPXux8WJ7WidoeaRudwbi5s5LeZ0D1Sw/pN1J4I3zneZ3F
eskvmSMuNmiWgXM71PinyMjLuqjLO52bvyf8CuYmndmhowzSV5UG8KkmoQN0y3Uf
+XEGLVuqM3dS4qZfXTGjruIjwVydGt0gY0omHokkMhHLb0N0WWaK4xN8EXtKzrOT
e27LG9byXPiaGJohMMXi93rw0uZ9w1IixduxInWKEBpRAn3rAtWvPBJPnn0M2Jy9
LrWunRzdF4PQ8k20YKdGnHx9DGv+7YfhHDTJmeYtoUXeQRNPIsogUv/gGI4zQy0K
HBRLUE3DU23mckueQyOnEA==

`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype="base64", line_length=64, bytes=3968)
`pragma protect data_block
aXGEOydeS5I+g0Yfv5+4dBlxKdFedb7019G2/J+a9I2ZSZHCJExKmpDDXKEZWAR2
kCkGdvundOQ76+pbp1yxNa+GJsEL0OSnSkelRKbh2DgF7a4s82TuEJoSM41TXmV7
XLP/zUitnuMJZiCcJax35MuBdjHzENpXVQ9NIgezPL+h6cvBMZkoTscFlgMF3AI6
tmyx4xAsrVVLkeDxK9WIfZLpEXAeg6MCHqurszuOGBFYLCh6vNPKRCHa9y03fQR5
Zuz5M3euYBp4uRiZKe1o8YdEnH40Rc/tTBfH2249XhHIg+eptRGuwrM11CEw1Qp9
e6J4GkYK/oPnmkEUTajyq3i0ko0/9VzklkRabW3h40ico4FMDXzdUVBUVaEGsarc
yLumg3IILcBjLEPBUd4WTgoJSnFoSbFoesagj79uOOGAALwF3Aqqoa3T9AsKN6AZ
oa3v+WyweNENTLP352N6/nq5O5ILjgAaYIWAWJ5+iOiWzY3FfVPVj2beRD/WVPUT
tp7cBeZCUBE23Ev+yG890fw1Xv7J5RCvTBWnSi29/oxIOtxBfRxG2KtpmhOxGijC
+2w0lOZuwNl8P2WkbAfL8YYmhiD+3OJ1r5PyVq1Xo/NDsCzVnCwLIVeRSmY/1saL
sotKHud62TtP60CiZzemHJVxek1wttohwVgECEZT4G9oEupQbXHBOV5vUvRKCDdP
L//CGoc+aoicpyjkX4ofcNRA+w/7W18csTTTsO3OU+Gsw9nMuPm6lGMeWzxSB74x
FDJZctA/fYjhYQBMptW6qFtCDXZsm0nq2cUA5V/ACN4ZGvsM3BfFd+31CvN/0y7A
UbbXCuBZFkNro6zEJzbKTJYCrWY0hGJILiZFoiN3Uy+TT42ofCebz3FdKb/usWi/
Ko+UxxwNF+0mmob9dhfOVvB+/8LNLl3H7rT66+J6LboW64E7DhEKGCpQNZn1+knr
D0m7fUIILyOChIykUSkL5fipsY0brBi9fmyiLBbw7JzEGOQASK81JrObyzkLxvpp
6Au5dP7Iw57WH0ouKXyKXP2E9+gQOAn/AZj6whgUpBh+EZEND2oyBATVjwKxkcau
00zEFZmKfbrz5AHh506FzaPTs2r23au9qNl1KyfGetpBp+gE7DFAqE/LnocV1zot
4HieKOKpomJEe03jVxQm0oIRJUiKEYUSnT/xqi0tCfxPm1aE+wKnhkzF+hscA02y
wB5CojnMzuK3u/McppssoyZ3144r4ZoOp5ct9aDOHy4Wmoq4A+rLqM8GA0u1L8nH
fSvpvqNhoP1uCoNGX5Vpns6BeoW2Y2S9Nor/Y/vWM7wai3achpy1y9UUl/T7nDSB
HzjAtSnylIjpUxtRC2PxTQc1LSLg5LQm0ti//nz8d+cukM3lvq8RV0Vf71+deRiu
LCHkDIhQcEiFZPW2agmPCz0iyj0iDGuy/v1vxNzo5IBYIQ3oFvG4iM0At8OUYkfF
eFJ8ubVpAuIAVZHD+rLyFuS/0aPU7kha6wwuRsvyv7Nq+Psojd8oHK7K0uxGO9ps
oCgZvDo1q9pdrOwMdyblKIRBtrVCo4ZGZmXCVkVqqI3YCTAVv8ut3cvjfTpHQHX3
9OJSTlRjV2T68ZvswGDZeZxewdIA3MbihVYdaBMkyLz5NijQ2kCz6Da1QEuqg74z
fC4NqxqfV41BWBQ6p6CkcCz63ONa7pBVV60tV2dC7W1MiKBtz7YuNS1CZNWdYb7n
5KzLGVkyeCO3ErqaQqUmH+gXJKxe7KDEEx4wmcETTngkF744AJmFU+JXp8BPGIEe
OvfWfG1RwpT98iUXHQ7hlzeiPtw5Pq6rRok+Zo/UNAcr4RaLBkuTnDAWt0VlC4Wk
y1Qn2J2gFmUUTA8Mmdp8l7WtDH3w1/qCweTTPt9rwU1bgDxxzEKc8n6JqYtunw++
KEb8gTEnZ5yN/yLkreUChruFH6z1/SMZejlsQ83z6Jib5qZkf1z7ITlYxrEuLYrE
6teDOJgsKnUyPYqcKuGzrhPLbDHl6CK1b3YGDCMkqe34hZxEpso9Gj7lY70wD3Ek
GLLHUt8m968WlBR5st9exNzI0pXQNDkGTpRcJmD1Jii2pq9fTiTkfdFTwAL+Dgrr
bwhMdGR9IrWfN3WdgP+SPYkRs8k+zad5orPL0bCULyaS04NNw0ZkHSNFoZVRxl+l
Qj/5TACyZKF1anPeDx64fqv98txxWG/fXNIRikr86nZbb8uB7Uqfk7vpO4kRDsCv
ZogD99HWvNnto0Q7TM2WzLC8sGZr1Ix7/gJVA/qlK96BSUxpGw/fTp97ub68Wf8P
0QD9RGRuc7UyofSX6jyn2Pzp8C2I20W7PM+y5jHOIQHrmod9cSHrqYlm/qyJaHFG
PCBZ23zbTAhBNBYAOjrlJBMfRif/yneCQj7FVcvZhOF3xe6l4e1/SEi/xx6CiX1b
RvsCeB23QkEjZaH408PMOnvkzS1f5CuSN43Y2ct22kPpK58A3gKSCpHWlyyHGlBj
cFPTg5xtPz3EA891HctZtAdfo6/+jV0ob+bSCRGVFbqYrM5avXgRn3b136Qg1NEY
ZlkGvHbEuSyoDVsWMA5sVTcgSfWeW3XMhYe3+/yU4MiT6aKxYNIouw+xE2Ug139O
oz1/ujaFXeiCGmwzUaUhGeQ/SqaxwjmQYyfqbtgOAj+URgr0WdFv5X2qPtP3+qIj
b7kAh3zRPldOEGZR8pBUzJ6Q/QVX6T9Mfncznk7mGVUsj4EPc28OwMBSRYII1f8m
lhRN4lodNYqlb47s1o0HUZOaicgR9JHrwpjrYJv79raEjzrZIg1+UHs4eqcAVhOC
92vNm4cxjCwC9/Z92lIDl3FCOH4Jr/he9gcB4n5rxMsNBmtpI7IAaRYcgIx6SiEq
6ZPyr5Ya7SAkDL33d7zheES/5Qa2UAtgLUcd8c6oJv4yBrpkaLxfviFtGzMs2Q1e
6UXiCItAYWH1aSj07YabA2rWcRiQSivg1Iyq0YlGS70XrdXD9O+l0av1UiYElZ4C
VtQ9Bm63e8PwhEwgmXX8nG29737WY88KcGkJspNPfjNJ0fFqghiUcrAR/Pck5i4s
leA+jVGjiqod4lqzISbaBPCIAwsszBf0ul+rCvBCBZqwRBqQEdobtKmlkrzEFxLN
k9PcbovrMDxFj3ArjsbLH5/FtSenr/73T9op+huISbQ1gvya7eaONQ2dej9EEL2s
jPKdUkZH//piwJq09s6g4jhunVodHfa4vQYZ0dfpVp/c4/VUiwFLR6LtfK0iPX50
w/jc28ABgRKCk+B2aMCqdTat7W9g3O15sokQzYXS1bC9X/Td4rG09h9BAcm7KmPe
U8LKIMj1X0y6LMFWmeZAPb4vLjgs/noCTzBgloFKpK99mAH+HonFplGKpF92F/fF
DxL24FYsSh71r/Uf93Hif1JJpKmQyF+7WQ+ygq+ErQfXXfxTaOumRRF9rrU20+2M
5uqytbEuL9ChBJ4l+Rn7JFb9pcRz28xfjG5RMGbasCFQkXP9NNml0CYS7NNca39V
GEBuT8aTZM1ITT707yApC6cGxohvGavCbztgI43S0dXWg7TBRgAlZkg+L7gnay11
UBQM/z8JEKRGVMZHl0tB8799OtnVBTgjGPSFD60cp7WAnPwPNh/mMrn/SFuBBqRs
XAcnP3+K58VULk3WgIYprnQVsDYqkYuK/sk9NyxO52X53ENwUofvdU66yyUiBY+x
OsHiIld6M1gMQfiHvFYsFEplbPxA/nYcTlDxkWar/eAuL5XO3N1lKU6IKIF0Nrkj
GhBHd79wBU72RDW4c97DyXRJkmIhLR2wCaN1jS5+6fXwckaouttxO8rFQF0DEmWw
dZRyQSLiNV7Qz7v/Gga+VRU22hwqeyppK/TYijpo2wP5xDev7e69MaICik0ePKPp
/KiMSEX2NNTWJraweqPwPm1+4jojzjVPpaWEWdHtEwH3hp1c+MqRu2P+2QnvYdbG
Hm0VJ5GybQ9DqGLg5sdZyMFTVN4jGPI/qqiu97Pew4nrJqJN0uspERIiBPEXc7mb
khZL8BCzwOT7CKUDfD6ku42bEq2bVEq1LiLYHUgafZ0gL5M1jOa7gyvod/Lc4kZG
JwIn6KkPCPC1opEl3rrzVCobE+H7IwBkItLGUzFYRqQ4JcEs9lwhLIXA3+0MD7NT
9igPNA+19u72l0sUWI5VPb5tx4OuC371pTisrcKIs3acagGqXqro38WHTA/AXs0u
Lay6LE6J1qeUIUn1UIviopT53SOWJ/FQ+j130XQgQGr0FwnyJa0vZS8hDNx62o8Y
DjbgprN5sTeziqixLnuzw8Qe9e4szbRhvOA5qdk4izvwrUT2uwosV4Oaibdyk7Gn
wkDw65EoMx6qu+EFuEYIDHYoe6Fz3+IlDVbKao0ddcJMX2GE+QlNqiFym3NrQFVH
lfJ+2NhrYv9vUfYKbjaQHP606kpCnWIggkJBbXiEGlIQ7VWSnueKnwYrfObb/KLv
21cBoAjXMVA5+BYaaeIVmDpCstha3L6DHdq1aV0VhWGZAp5LdWFOXGx9RLceC4Ww
rOAk+k9Kh2+NBQeKLQO9E/j+AGoSI2SP0DDlUchn2KY+moDoFWg8AgSx66vo1Sdk
nXXyFykJ3HnkHqm8+31+KZnf6yGiPBTs6EPYcy49NMoxFh0yJmnlSwMrVUaC7ZP0
fenWqfWYUV4bQnY2mtlBCjRCtXUE4XCegnlPMleGFY45rL9WEZ0sOXgMvJ7dhcMx
EqMLW04qWEKjRUOIHwIV2BZ0e6RTQLGfXCR/0sKpOHPtBgc9iOqfOspPYdwOZB5j
Kd6KLaQRYJaOhy2qfm6RKwxlwn6b4UQc2lQe487JVJ/Kc0uBJ4VEfY7sCqVxjP+4
lP+jgDx6hWRR3Jlips4/RKRz10sW9gmnUDg3JS505RRUC1+EuTyiUBp9m6/wryXZ
lwkI63bBkOSGQhv4CV+kx2s+iy6Xx8pTZS/2f38UPQ1AhkVrxW5+0ku2doQAsGqo
qs4PC5rvexSXMHDEdZKc+iUMjMGylrO8TFw9mV3onBgB0BwAT99KbUGchZCFNwsX
CEo8GIOcFO7/gnu0TvgIuK061uIiUbduFNPAXesRiumOj9btkQpGdxSF15E4nOkP
hGBvNmSGabemQX4YwhASHAPkS41HBZLI1DYOcCliOx1nkW5Do1MAmXGNmqbJfX8p
TAZwnmF+lWWx9NBSz8ce2RKmC+ZJc3RGVM6hxlIlNGrWTL31GKfNSkeE7abFjKHR
wnI5XJKMzjzuPpx4n87FLB3Nj7TiK4fTDQrNa0UOOTI=

`pragma protect end_protected
endmodule

