`timescale 1ps/1ps
module RAM40_16K ( RDATA, RCLK, RCLKE, RE, RADDR, WCLK, WCLKE, WE, WADDR, MASK, WDATA ); 

output	[15:0]	RDATA;  
input         	RCLK;   
input           RCLKE; 
input           RE; 
input	[12:0]  RADDR; 
input           WCLK; 
input           WCLKE; 
input           WE; 
input 	[12:0]  WADDR; 
input 	[15:0]  MASK; 
input 	[15:0]	WDATA; 


parameter WRITE_MODE = 0;    // Configure Write Port as 1024x16 (0)/ 20148x8 (1)/ 4096x4 (2)/ 8192x2 (3)     
parameter READ_MODE  = 0;    // Configure Read  Port as 1024x16 (0)/ 20148x8 (1)/ 4096x4 (2)/ 8192x2 (3)

parameter INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

parameter INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
parameter INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;  
 

assign (weak0, weak1) MASK = 16'b0;

wire [15:0] RD;
wire [15:0] WD;
wire [15:0] MASK_RAM;

reg [12:10] RADDR_reg;
always @(posedge RCLK) begin
	RADDR_reg[12:10] <= RADDR[12:10];
end

read_data_decoder read_decoder_inst (
	.di(RD),
	.ai(RADDR_reg[12:10]),
	.do(RDATA)
);
defparam read_decoder_inst.READ_MODE = READ_MODE;

write_data_decoder write_decoder_inst (
	.di(WDATA),
	.do(WD)
);
defparam write_decoder_inst.WRITE_MODE = WRITE_MODE;

mask_decoder mask_decoder_inst(
	.mi(MASK),
	.ai(WADDR[12:10]),
	.mo(MASK_RAM)
);
defparam mask_decoder_inst.WRITE_MODE = WRITE_MODE;

RAM16K ram_inst (
	.RDATA(RD),
	.RCLK(RCLK),
	.RCLKE(RCLKE),
	.RE(RE),
	.RADDR(RADDR[9:0]),
	.WCLK(WCLK),
	.WCLKE(WCLKE),
	.WE(WE),
	.WADDR(WADDR[9:0]),
	.MASK(MASK_RAM),
	.WDATA(WD));

defparam ram_inst.INIT_0 = INIT_0;
defparam ram_inst.INIT_1 = INIT_1;
defparam ram_inst.INIT_2 = INIT_2;
defparam ram_inst.INIT_3 = INIT_3;
defparam ram_inst.INIT_4 = INIT_4;
defparam ram_inst.INIT_5 = INIT_5;
defparam ram_inst.INIT_6 = INIT_6;
defparam ram_inst.INIT_7 = INIT_7;
defparam ram_inst.INIT_8 = INIT_8;
defparam ram_inst.INIT_9 = INIT_9;
defparam ram_inst.INIT_A = INIT_A;
defparam ram_inst.INIT_B = INIT_B;
defparam ram_inst.INIT_C = INIT_C;
defparam ram_inst.INIT_D = INIT_D;
defparam ram_inst.INIT_E = INIT_E;
defparam ram_inst.INIT_F = INIT_F;

defparam ram_inst.INIT_10 = INIT_10;
defparam ram_inst.INIT_11 = INIT_11;
defparam ram_inst.INIT_12 = INIT_12;
defparam ram_inst.INIT_13 = INIT_13;
defparam ram_inst.INIT_14 = INIT_14;
defparam ram_inst.INIT_15 = INIT_15;
defparam ram_inst.INIT_16 = INIT_16;
defparam ram_inst.INIT_17 = INIT_17;
defparam ram_inst.INIT_18 = INIT_18;
defparam ram_inst.INIT_19 = INIT_19;
defparam ram_inst.INIT_1A = INIT_1A;
defparam ram_inst.INIT_1B = INIT_1B;
defparam ram_inst.INIT_1C = INIT_1C;
defparam ram_inst.INIT_1D = INIT_1D;
defparam ram_inst.INIT_1E = INIT_1E;
defparam ram_inst.INIT_1F = INIT_1F;

defparam ram_inst.INIT_20 = INIT_20;
defparam ram_inst.INIT_21 = INIT_21;
defparam ram_inst.INIT_22 = INIT_22;
defparam ram_inst.INIT_23 = INIT_23;
defparam ram_inst.INIT_24 = INIT_24;
defparam ram_inst.INIT_25 = INIT_25;
defparam ram_inst.INIT_26 = INIT_26;
defparam ram_inst.INIT_27 = INIT_27;
defparam ram_inst.INIT_28 = INIT_28;
defparam ram_inst.INIT_29 = INIT_29;
defparam ram_inst.INIT_2A = INIT_2A;
defparam ram_inst.INIT_2B = INIT_2B;
defparam ram_inst.INIT_2C = INIT_2C;
defparam ram_inst.INIT_2D = INIT_2D;
defparam ram_inst.INIT_2E = INIT_2E;
defparam ram_inst.INIT_2F = INIT_2F;

defparam ram_inst.INIT_30 = INIT_30;
defparam ram_inst.INIT_31 = INIT_31;
defparam ram_inst.INIT_32 = INIT_32;
defparam ram_inst.INIT_33 = INIT_33;
defparam ram_inst.INIT_34 = INIT_34;
defparam ram_inst.INIT_35 = INIT_35;
defparam ram_inst.INIT_36 = INIT_36;
defparam ram_inst.INIT_37 = INIT_37;
defparam ram_inst.INIT_38 = INIT_38;
defparam ram_inst.INIT_39 = INIT_39;
defparam ram_inst.INIT_3A = INIT_3A;
defparam ram_inst.INIT_3B = INIT_3B;
defparam ram_inst.INIT_3C = INIT_3C;
defparam ram_inst.INIT_3D = INIT_3D;
defparam ram_inst.INIT_3E = INIT_3E;
defparam ram_inst.INIT_3F = INIT_3F;


endmodule // RAM40_16K;
