`timescale 1ps/1ps
module IR_IP(
// *** Input to UUT ***
 input            IRIN,
 input            ADRI3,
 input            ADRI2,
 input            ADRI1,
 input            ADRI0,
 input            CSI,
 input            DENI,
 input            EXE,
 input            LEARN,
 input            RST,
 input            WEI,
 input  		  CLKI,
// *** Outputs from UUT ***
 output            IROUT,
 output            BUSY,
 output            DRDY,
 output            ERR,
 output            RDATA0,
 output            RDATA1,
 output            RDATA2,
 output            RDATA3,
 output            RDATA4,
 output            RDATA5,
 output            RDATA6,
 output            RDATA7,


 input            WDATA0,
 input            WDATA1,
 input            WDATA2,
 input            WDATA3,
 input            WDATA4,
 input            WDATA5,
 input            WDATA6,
 input            WDATA7
 );

IR_IP_CORE inst (
			 .CLKI(CLKI),
             .IRIN(IRIN),
             .ADRI3(ADRI3),
             .ADRI2(ADRI2),
             .ADRI1(ADRI1),
             .ADRI0(ADRI0),
             .CSI(CSI),
             .DENI(DENI),
             .EXE(EXE),
             .LEARN(LEARN),
             .RST(RST),
             .WEI(WEI),
             .IROUT(IROUT),
             .BUSY(BUSY),
             .DRDY(DRDY),
             .ERR(ERR),
             .RDATA0(RDATA0),
             .RDATA1(RDATA1),
             .RDATA2(RDATA2),
             .RDATA3(RDATA3),
             .RDATA4(RDATA4),
             .RDATA5(RDATA5),
             .RDATA6(RDATA6),
             .RDATA7(RDATA7),
             .WDATA0(WDATA0),
             .WDATA1(WDATA1),
             .WDATA2(WDATA2),
             .WDATA3(WDATA3),
             .WDATA4(WDATA4),
             .WDATA5(WDATA5),
             .WDATA6(WDATA6),
             .WDATA7(WDATA7)
);
 endmodule
