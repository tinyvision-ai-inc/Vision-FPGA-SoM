`timescale 1ns/1ns
module VHI ( Z );
    output Z ;
  supply1 VSS;
  buf (Z , VSS);
endmodule
