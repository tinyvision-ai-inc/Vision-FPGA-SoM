`timescale 10ps/1ps
module LocalMux(I, O);
input I;
output O;


	assign O = I;
endmodule
