`timescale 10ps/1ps
module CEMux(I, O);
input I;
output O;

	assign O = I;


endmodule
