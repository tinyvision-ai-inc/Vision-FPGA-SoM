`timescale 1ps/1ps
module GND (Y);

    output Y;
supply0 Y ;
endmodule
