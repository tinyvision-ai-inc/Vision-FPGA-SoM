`timescale 10ps/1ps
module Odrv12(I, O);
input I;
output O;

	assign O = I;
	

endmodule
