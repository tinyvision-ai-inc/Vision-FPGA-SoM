`timescale 10ps/1ps
module Odrv4(I, O);
input I;
output O;

	assign O = I;


endmodule
