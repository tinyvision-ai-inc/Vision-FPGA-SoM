`timescale 10ps/1ps
module Span4Mux_s2_h(I, O);
input I;
output O;

	assign O = I;
	

endmodule
