`timescale 1ns / 10ps 
module esd_btbdiodes ( vssx );

  input vssx;
endmodule
