`timescale 1ps/1ps
module BARCODE_DRV   (
	CURREN,
	BARCODEEN,
	BARCODEPWM,
	BARCODE
);

parameter BARCODE_CURRENT = "0b0000";
parameter CURRENT_MODE = "0b0";

	input CURREN,	BARCODEEN, 	BARCODEPWM; 
	output 	BARCODE; 

 BARCODE_DRV_CORE #(.BARCODE_CURRENT(BARCODE_CURRENT),.CURRENT_MODE(CURRENT_MODE))
inst
 (
	.CURREN(CURREN),
	.BARCODEEN(BARCODEEN),
	.BARCODEPWM(BARCODEPWM),
	.BARCODE(BARCODE)
);

endmodule
