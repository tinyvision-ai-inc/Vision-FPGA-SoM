`timescale 1ps/1ps
module GB (	
GLOBAL_BUFFER_OUTPUT,
USER_SIGNAL_TO_GLOBAL_BUFFER);

input USER_SIGNAL_TO_GLOBAL_BUFFER;			
output GLOBAL_BUFFER_OUTPUT;	

assign GLOBAL_BUFFER_OUTPUT = USER_SIGNAL_TO_GLOBAL_BUFFER;



endmodule	//GB
