`timescale 10ps/1ps
module CascadeMux(I, O);
input I;
output O;

assign O = I;


endmodule
